-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 13 2023 19:34:34

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "test" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of test
entity test is
port (
    LED4 : out std_logic;
    LED2 : out std_logic;
    LED5 : out std_logic;
    LED3 : out std_logic;
    LED1 : out std_logic);
end test;

-- Architecture of test
-- View name is \INTERFACE\
architecture \INTERFACE\ of test is

signal \N__9920\ : std_logic;
signal \N__9919\ : std_logic;
signal \N__9918\ : std_logic;
signal \N__9911\ : std_logic;
signal \N__9910\ : std_logic;
signal \N__9909\ : std_logic;
signal \N__9902\ : std_logic;
signal \N__9901\ : std_logic;
signal \N__9900\ : std_logic;
signal \N__9893\ : std_logic;
signal \N__9892\ : std_logic;
signal \N__9891\ : std_logic;
signal \N__9884\ : std_logic;
signal \N__9883\ : std_logic;
signal \N__9882\ : std_logic;
signal \N__9865\ : std_logic;
signal \N__9862\ : std_logic;
signal \N__9859\ : std_logic;
signal \N__9856\ : std_logic;
signal \N__9853\ : std_logic;
signal \N__9852\ : std_logic;
signal \N__9851\ : std_logic;
signal \N__9850\ : std_logic;
signal \N__9847\ : std_logic;
signal \N__9844\ : std_logic;
signal \N__9841\ : std_logic;
signal \N__9840\ : std_logic;
signal \N__9837\ : std_logic;
signal \N__9836\ : std_logic;
signal \N__9829\ : std_logic;
signal \N__9826\ : std_logic;
signal \N__9823\ : std_logic;
signal \N__9820\ : std_logic;
signal \N__9815\ : std_logic;
signal \N__9808\ : std_logic;
signal \N__9805\ : std_logic;
signal \N__9804\ : std_logic;
signal \N__9803\ : std_logic;
signal \N__9802\ : std_logic;
signal \N__9799\ : std_logic;
signal \N__9796\ : std_logic;
signal \N__9793\ : std_logic;
signal \N__9790\ : std_logic;
signal \N__9785\ : std_logic;
signal \N__9782\ : std_logic;
signal \N__9779\ : std_logic;
signal \N__9772\ : std_logic;
signal \N__9771\ : std_logic;
signal \N__9768\ : std_logic;
signal \N__9767\ : std_logic;
signal \N__9764\ : std_logic;
signal \N__9763\ : std_logic;
signal \N__9760\ : std_logic;
signal \N__9757\ : std_logic;
signal \N__9754\ : std_logic;
signal \N__9751\ : std_logic;
signal \N__9748\ : std_logic;
signal \N__9743\ : std_logic;
signal \N__9740\ : std_logic;
signal \N__9739\ : std_logic;
signal \N__9736\ : std_logic;
signal \N__9733\ : std_logic;
signal \N__9730\ : std_logic;
signal \N__9727\ : std_logic;
signal \N__9718\ : std_logic;
signal \N__9715\ : std_logic;
signal \N__9714\ : std_logic;
signal \N__9713\ : std_logic;
signal \N__9712\ : std_logic;
signal \N__9711\ : std_logic;
signal \N__9708\ : std_logic;
signal \N__9705\ : std_logic;
signal \N__9702\ : std_logic;
signal \N__9697\ : std_logic;
signal \N__9692\ : std_logic;
signal \N__9687\ : std_logic;
signal \N__9684\ : std_logic;
signal \N__9681\ : std_logic;
signal \N__9676\ : std_logic;
signal \N__9675\ : std_logic;
signal \N__9672\ : std_logic;
signal \N__9671\ : std_logic;
signal \N__9670\ : std_logic;
signal \N__9667\ : std_logic;
signal \N__9666\ : std_logic;
signal \N__9665\ : std_logic;
signal \N__9656\ : std_logic;
signal \N__9655\ : std_logic;
signal \N__9654\ : std_logic;
signal \N__9653\ : std_logic;
signal \N__9652\ : std_logic;
signal \N__9651\ : std_logic;
signal \N__9650\ : std_logic;
signal \N__9645\ : std_logic;
signal \N__9642\ : std_logic;
signal \N__9637\ : std_logic;
signal \N__9632\ : std_logic;
signal \N__9629\ : std_logic;
signal \N__9626\ : std_logic;
signal \N__9613\ : std_logic;
signal \N__9612\ : std_logic;
signal \N__9611\ : std_logic;
signal \N__9610\ : std_logic;
signal \N__9609\ : std_logic;
signal \N__9608\ : std_logic;
signal \N__9607\ : std_logic;
signal \N__9604\ : std_logic;
signal \N__9601\ : std_logic;
signal \N__9600\ : std_logic;
signal \N__9597\ : std_logic;
signal \N__9594\ : std_logic;
signal \N__9591\ : std_logic;
signal \N__9590\ : std_logic;
signal \N__9589\ : std_logic;
signal \N__9586\ : std_logic;
signal \N__9577\ : std_logic;
signal \N__9572\ : std_logic;
signal \N__9571\ : std_logic;
signal \N__9566\ : std_logic;
signal \N__9561\ : std_logic;
signal \N__9556\ : std_logic;
signal \N__9553\ : std_logic;
signal \N__9544\ : std_logic;
signal \N__9543\ : std_logic;
signal \N__9540\ : std_logic;
signal \N__9539\ : std_logic;
signal \N__9536\ : std_logic;
signal \N__9535\ : std_logic;
signal \N__9530\ : std_logic;
signal \N__9527\ : std_logic;
signal \N__9526\ : std_logic;
signal \N__9525\ : std_logic;
signal \N__9524\ : std_logic;
signal \N__9523\ : std_logic;
signal \N__9522\ : std_logic;
signal \N__9521\ : std_logic;
signal \N__9520\ : std_logic;
signal \N__9517\ : std_logic;
signal \N__9512\ : std_logic;
signal \N__9509\ : std_logic;
signal \N__9500\ : std_logic;
signal \N__9495\ : std_logic;
signal \N__9490\ : std_logic;
signal \N__9481\ : std_logic;
signal \N__9478\ : std_logic;
signal \N__9475\ : std_logic;
signal \N__9472\ : std_logic;
signal \N__9469\ : std_logic;
signal \N__9468\ : std_logic;
signal \N__9465\ : std_logic;
signal \N__9464\ : std_logic;
signal \N__9461\ : std_logic;
signal \N__9460\ : std_logic;
signal \N__9459\ : std_logic;
signal \N__9458\ : std_logic;
signal \N__9455\ : std_logic;
signal \N__9452\ : std_logic;
signal \N__9449\ : std_logic;
signal \N__9446\ : std_logic;
signal \N__9441\ : std_logic;
signal \N__9436\ : std_logic;
signal \N__9427\ : std_logic;
signal \N__9424\ : std_logic;
signal \N__9421\ : std_logic;
signal \N__9420\ : std_logic;
signal \N__9419\ : std_logic;
signal \N__9416\ : std_logic;
signal \N__9413\ : std_logic;
signal \N__9410\ : std_logic;
signal \N__9403\ : std_logic;
signal \N__9402\ : std_logic;
signal \N__9401\ : std_logic;
signal \N__9400\ : std_logic;
signal \N__9397\ : std_logic;
signal \N__9396\ : std_logic;
signal \N__9395\ : std_logic;
signal \N__9394\ : std_logic;
signal \N__9393\ : std_logic;
signal \N__9390\ : std_logic;
signal \N__9387\ : std_logic;
signal \N__9384\ : std_logic;
signal \N__9381\ : std_logic;
signal \N__9378\ : std_logic;
signal \N__9373\ : std_logic;
signal \N__9370\ : std_logic;
signal \N__9367\ : std_logic;
signal \N__9364\ : std_logic;
signal \N__9363\ : std_logic;
signal \N__9362\ : std_logic;
signal \N__9357\ : std_logic;
signal \N__9356\ : std_logic;
signal \N__9353\ : std_logic;
signal \N__9350\ : std_logic;
signal \N__9345\ : std_logic;
signal \N__9342\ : std_logic;
signal \N__9337\ : std_logic;
signal \N__9334\ : std_logic;
signal \N__9331\ : std_logic;
signal \N__9324\ : std_logic;
signal \N__9313\ : std_logic;
signal \N__9310\ : std_logic;
signal \N__9309\ : std_logic;
signal \N__9306\ : std_logic;
signal \N__9303\ : std_logic;
signal \N__9298\ : std_logic;
signal \N__9297\ : std_logic;
signal \N__9294\ : std_logic;
signal \N__9291\ : std_logic;
signal \N__9286\ : std_logic;
signal \N__9283\ : std_logic;
signal \N__9280\ : std_logic;
signal \N__9279\ : std_logic;
signal \N__9278\ : std_logic;
signal \N__9275\ : std_logic;
signal \N__9270\ : std_logic;
signal \N__9265\ : std_logic;
signal \N__9262\ : std_logic;
signal \N__9259\ : std_logic;
signal \N__9258\ : std_logic;
signal \N__9255\ : std_logic;
signal \N__9252\ : std_logic;
signal \N__9247\ : std_logic;
signal \N__9244\ : std_logic;
signal \N__9241\ : std_logic;
signal \N__9240\ : std_logic;
signal \N__9239\ : std_logic;
signal \N__9236\ : std_logic;
signal \N__9233\ : std_logic;
signal \N__9230\ : std_logic;
signal \N__9227\ : std_logic;
signal \N__9224\ : std_logic;
signal \N__9221\ : std_logic;
signal \N__9220\ : std_logic;
signal \N__9217\ : std_logic;
signal \N__9212\ : std_logic;
signal \N__9209\ : std_logic;
signal \N__9206\ : std_logic;
signal \N__9201\ : std_logic;
signal \N__9196\ : std_logic;
signal \N__9195\ : std_logic;
signal \N__9194\ : std_logic;
signal \N__9191\ : std_logic;
signal \N__9188\ : std_logic;
signal \N__9185\ : std_logic;
signal \N__9182\ : std_logic;
signal \N__9179\ : std_logic;
signal \N__9176\ : std_logic;
signal \N__9175\ : std_logic;
signal \N__9172\ : std_logic;
signal \N__9169\ : std_logic;
signal \N__9166\ : std_logic;
signal \N__9163\ : std_logic;
signal \N__9158\ : std_logic;
signal \N__9155\ : std_logic;
signal \N__9152\ : std_logic;
signal \N__9147\ : std_logic;
signal \N__9144\ : std_logic;
signal \N__9139\ : std_logic;
signal \N__9138\ : std_logic;
signal \N__9137\ : std_logic;
signal \N__9134\ : std_logic;
signal \N__9133\ : std_logic;
signal \N__9130\ : std_logic;
signal \N__9127\ : std_logic;
signal \N__9124\ : std_logic;
signal \N__9123\ : std_logic;
signal \N__9120\ : std_logic;
signal \N__9117\ : std_logic;
signal \N__9114\ : std_logic;
signal \N__9111\ : std_logic;
signal \N__9110\ : std_logic;
signal \N__9107\ : std_logic;
signal \N__9104\ : std_logic;
signal \N__9101\ : std_logic;
signal \N__9098\ : std_logic;
signal \N__9095\ : std_logic;
signal \N__9092\ : std_logic;
signal \N__9079\ : std_logic;
signal \N__9078\ : std_logic;
signal \N__9077\ : std_logic;
signal \N__9076\ : std_logic;
signal \N__9075\ : std_logic;
signal \N__9074\ : std_logic;
signal \N__9073\ : std_logic;
signal \N__9072\ : std_logic;
signal \N__9071\ : std_logic;
signal \N__9068\ : std_logic;
signal \N__9065\ : std_logic;
signal \N__9058\ : std_logic;
signal \N__9055\ : std_logic;
signal \N__9054\ : std_logic;
signal \N__9053\ : std_logic;
signal \N__9050\ : std_logic;
signal \N__9047\ : std_logic;
signal \N__9046\ : std_logic;
signal \N__9045\ : std_logic;
signal \N__9044\ : std_logic;
signal \N__9043\ : std_logic;
signal \N__9042\ : std_logic;
signal \N__9039\ : std_logic;
signal \N__9038\ : std_logic;
signal \N__9037\ : std_logic;
signal \N__9034\ : std_logic;
signal \N__9033\ : std_logic;
signal \N__9032\ : std_logic;
signal \N__9029\ : std_logic;
signal \N__9026\ : std_logic;
signal \N__9023\ : std_logic;
signal \N__9020\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9012\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9006\ : std_logic;
signal \N__9005\ : std_logic;
signal \N__9002\ : std_logic;
signal \N__8995\ : std_logic;
signal \N__8992\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8986\ : std_logic;
signal \N__8985\ : std_logic;
signal \N__8984\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8978\ : std_logic;
signal \N__8977\ : std_logic;
signal \N__8976\ : std_logic;
signal \N__8975\ : std_logic;
signal \N__8974\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8968\ : std_logic;
signal \N__8961\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8951\ : std_logic;
signal \N__8948\ : std_logic;
signal \N__8941\ : std_logic;
signal \N__8938\ : std_logic;
signal \N__8935\ : std_logic;
signal \N__8932\ : std_logic;
signal \N__8929\ : std_logic;
signal \N__8924\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8917\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8905\ : std_logic;
signal \N__8902\ : std_logic;
signal \N__8897\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8880\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8851\ : std_logic;
signal \N__8850\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8847\ : std_logic;
signal \N__8846\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8844\ : std_logic;
signal \N__8843\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8828\ : std_logic;
signal \N__8827\ : std_logic;
signal \N__8822\ : std_logic;
signal \N__8817\ : std_logic;
signal \N__8812\ : std_logic;
signal \N__8809\ : std_logic;
signal \N__8800\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8793\ : std_logic;
signal \N__8790\ : std_logic;
signal \N__8787\ : std_logic;
signal \N__8784\ : std_logic;
signal \N__8781\ : std_logic;
signal \N__8778\ : std_logic;
signal \N__8773\ : std_logic;
signal \N__8770\ : std_logic;
signal \N__8769\ : std_logic;
signal \N__8768\ : std_logic;
signal \N__8767\ : std_logic;
signal \N__8766\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8762\ : std_logic;
signal \N__8761\ : std_logic;
signal \N__8758\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8753\ : std_logic;
signal \N__8750\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8744\ : std_logic;
signal \N__8741\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8730\ : std_logic;
signal \N__8727\ : std_logic;
signal \N__8724\ : std_logic;
signal \N__8721\ : std_logic;
signal \N__8718\ : std_logic;
signal \N__8717\ : std_logic;
signal \N__8716\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8710\ : std_logic;
signal \N__8707\ : std_logic;
signal \N__8704\ : std_logic;
signal \N__8695\ : std_logic;
signal \N__8692\ : std_logic;
signal \N__8689\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8670\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8658\ : std_logic;
signal \N__8657\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8643\ : std_logic;
signal \N__8638\ : std_logic;
signal \N__8635\ : std_logic;
signal \N__8634\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8627\ : std_logic;
signal \N__8624\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8616\ : std_logic;
signal \N__8611\ : std_logic;
signal \N__8602\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8598\ : std_logic;
signal \N__8597\ : std_logic;
signal \N__8594\ : std_logic;
signal \N__8591\ : std_logic;
signal \N__8586\ : std_logic;
signal \N__8581\ : std_logic;
signal \N__8580\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8578\ : std_logic;
signal \N__8577\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8575\ : std_logic;
signal \N__8574\ : std_logic;
signal \N__8569\ : std_logic;
signal \N__8566\ : std_logic;
signal \N__8559\ : std_logic;
signal \N__8556\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8546\ : std_logic;
signal \N__8541\ : std_logic;
signal \N__8536\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8525\ : std_logic;
signal \N__8522\ : std_logic;
signal \N__8515\ : std_logic;
signal \N__8510\ : std_logic;
signal \N__8503\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8497\ : std_logic;
signal \N__8496\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8492\ : std_logic;
signal \N__8489\ : std_logic;
signal \N__8488\ : std_logic;
signal \N__8485\ : std_logic;
signal \N__8482\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8477\ : std_logic;
signal \N__8474\ : std_logic;
signal \N__8471\ : std_logic;
signal \N__8466\ : std_logic;
signal \N__8465\ : std_logic;
signal \N__8464\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8455\ : std_logic;
signal \N__8450\ : std_logic;
signal \N__8445\ : std_logic;
signal \N__8442\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8430\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8423\ : std_logic;
signal \N__8420\ : std_logic;
signal \N__8417\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8405\ : std_logic;
signal \N__8404\ : std_logic;
signal \N__8401\ : std_logic;
signal \N__8398\ : std_logic;
signal \N__8393\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8385\ : std_logic;
signal \N__8384\ : std_logic;
signal \N__8383\ : std_logic;
signal \N__8382\ : std_logic;
signal \N__8379\ : std_logic;
signal \N__8376\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8372\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8366\ : std_logic;
signal \N__8361\ : std_logic;
signal \N__8360\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8329\ : std_logic;
signal \N__8324\ : std_logic;
signal \N__8321\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8305\ : std_logic;
signal \N__8302\ : std_logic;
signal \N__8301\ : std_logic;
signal \N__8298\ : std_logic;
signal \N__8295\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8287\ : std_logic;
signal \N__8286\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8282\ : std_logic;
signal \N__8281\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8278\ : std_logic;
signal \N__8275\ : std_logic;
signal \N__8274\ : std_logic;
signal \N__8273\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8271\ : std_logic;
signal \N__8268\ : std_logic;
signal \N__8265\ : std_logic;
signal \N__8262\ : std_logic;
signal \N__8261\ : std_logic;
signal \N__8260\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8250\ : std_logic;
signal \N__8247\ : std_logic;
signal \N__8242\ : std_logic;
signal \N__8239\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8226\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8218\ : std_logic;
signal \N__8215\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8205\ : std_logic;
signal \N__8200\ : std_logic;
signal \N__8197\ : std_logic;
signal \N__8194\ : std_logic;
signal \N__8191\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8178\ : std_logic;
signal \N__8175\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8157\ : std_logic;
signal \N__8154\ : std_logic;
signal \N__8151\ : std_logic;
signal \N__8148\ : std_logic;
signal \N__8145\ : std_logic;
signal \N__8140\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8128\ : std_logic;
signal \N__8125\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8112\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8108\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8099\ : std_logic;
signal \N__8098\ : std_logic;
signal \N__8095\ : std_logic;
signal \N__8092\ : std_logic;
signal \N__8089\ : std_logic;
signal \N__8086\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8074\ : std_logic;
signal \N__8073\ : std_logic;
signal \N__8070\ : std_logic;
signal \N__8067\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8063\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8050\ : std_logic;
signal \N__8047\ : std_logic;
signal \N__8044\ : std_logic;
signal \N__8043\ : std_logic;
signal \N__8038\ : std_logic;
signal \N__8035\ : std_logic;
signal \N__8032\ : std_logic;
signal \N__8031\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8027\ : std_logic;
signal \N__8024\ : std_logic;
signal \N__8023\ : std_logic;
signal \N__8020\ : std_logic;
signal \N__8017\ : std_logic;
signal \N__8014\ : std_logic;
signal \N__8011\ : std_logic;
signal \N__8008\ : std_logic;
signal \N__8005\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7987\ : std_logic;
signal \N__7986\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7979\ : std_logic;
signal \N__7976\ : std_logic;
signal \N__7975\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7966\ : std_logic;
signal \N__7965\ : std_logic;
signal \N__7962\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7954\ : std_logic;
signal \N__7949\ : std_logic;
signal \N__7946\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7935\ : std_logic;
signal \N__7934\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7930\ : std_logic;
signal \N__7929\ : std_logic;
signal \N__7926\ : std_logic;
signal \N__7921\ : std_logic;
signal \N__7918\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7912\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7899\ : std_logic;
signal \N__7894\ : std_logic;
signal \N__7893\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7880\ : std_logic;
signal \N__7877\ : std_logic;
signal \N__7874\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7872\ : std_logic;
signal \N__7869\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7859\ : std_logic;
signal \N__7852\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7846\ : std_logic;
signal \N__7843\ : std_logic;
signal \N__7840\ : std_logic;
signal \N__7837\ : std_logic;
signal \N__7836\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7827\ : std_logic;
signal \N__7824\ : std_logic;
signal \N__7821\ : std_logic;
signal \N__7818\ : std_logic;
signal \N__7813\ : std_logic;
signal \N__7810\ : std_logic;
signal \N__7807\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7791\ : std_logic;
signal \N__7786\ : std_logic;
signal \N__7783\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7780\ : std_logic;
signal \N__7779\ : std_logic;
signal \N__7776\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7765\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7763\ : std_logic;
signal \N__7762\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7760\ : std_logic;
signal \N__7759\ : std_logic;
signal \N__7758\ : std_logic;
signal \N__7755\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7739\ : std_logic;
signal \N__7736\ : std_logic;
signal \N__7733\ : std_logic;
signal \N__7728\ : std_logic;
signal \N__7725\ : std_logic;
signal \N__7722\ : std_logic;
signal \N__7715\ : std_logic;
signal \N__7708\ : std_logic;
signal \N__7699\ : std_logic;
signal \N__7696\ : std_logic;
signal \N__7693\ : std_logic;
signal \N__7692\ : std_logic;
signal \N__7689\ : std_logic;
signal \N__7688\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7684\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7677\ : std_logic;
signal \N__7674\ : std_logic;
signal \N__7671\ : std_logic;
signal \N__7668\ : std_logic;
signal \N__7665\ : std_logic;
signal \N__7662\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7652\ : std_logic;
signal \N__7645\ : std_logic;
signal \N__7644\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7640\ : std_logic;
signal \N__7637\ : std_logic;
signal \N__7636\ : std_logic;
signal \N__7633\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7623\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7617\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7596\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7589\ : std_logic;
signal \N__7586\ : std_logic;
signal \N__7583\ : std_logic;
signal \N__7580\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7571\ : std_logic;
signal \N__7568\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7562\ : std_logic;
signal \N__7559\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7549\ : std_logic;
signal \N__7548\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7538\ : std_logic;
signal \N__7535\ : std_logic;
signal \N__7532\ : std_logic;
signal \N__7529\ : std_logic;
signal \N__7526\ : std_logic;
signal \N__7523\ : std_logic;
signal \N__7516\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7514\ : std_logic;
signal \N__7511\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7504\ : std_logic;
signal \N__7503\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7497\ : std_logic;
signal \N__7494\ : std_logic;
signal \N__7491\ : std_logic;
signal \N__7488\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7482\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7450\ : std_logic;
signal \N__7447\ : std_logic;
signal \N__7444\ : std_logic;
signal \N__7439\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7429\ : std_logic;
signal \N__7428\ : std_logic;
signal \N__7425\ : std_logic;
signal \N__7422\ : std_logic;
signal \N__7421\ : std_logic;
signal \N__7420\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7418\ : std_logic;
signal \N__7417\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7415\ : std_logic;
signal \N__7414\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7407\ : std_logic;
signal \N__7406\ : std_logic;
signal \N__7405\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7403\ : std_logic;
signal \N__7402\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7392\ : std_logic;
signal \N__7387\ : std_logic;
signal \N__7386\ : std_logic;
signal \N__7383\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7372\ : std_logic;
signal \N__7369\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7360\ : std_logic;
signal \N__7357\ : std_logic;
signal \N__7354\ : std_logic;
signal \N__7351\ : std_logic;
signal \N__7348\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7329\ : std_logic;
signal \N__7328\ : std_logic;
signal \N__7327\ : std_logic;
signal \N__7324\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7285\ : std_logic;
signal \N__7278\ : std_logic;
signal \N__7269\ : std_logic;
signal \N__7258\ : std_logic;
signal \N__7255\ : std_logic;
signal \N__7254\ : std_logic;
signal \N__7251\ : std_logic;
signal \N__7248\ : std_logic;
signal \N__7247\ : std_logic;
signal \N__7244\ : std_logic;
signal \N__7239\ : std_logic;
signal \N__7238\ : std_logic;
signal \N__7237\ : std_logic;
signal \N__7234\ : std_logic;
signal \N__7231\ : std_logic;
signal \N__7228\ : std_logic;
signal \N__7225\ : std_logic;
signal \N__7222\ : std_logic;
signal \N__7217\ : std_logic;
signal \N__7210\ : std_logic;
signal \N__7209\ : std_logic;
signal \N__7206\ : std_logic;
signal \N__7203\ : std_logic;
signal \N__7200\ : std_logic;
signal \N__7197\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7189\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7185\ : std_logic;
signal \N__7182\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7171\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7164\ : std_logic;
signal \N__7163\ : std_logic;
signal \N__7160\ : std_logic;
signal \N__7157\ : std_logic;
signal \N__7154\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7141\ : std_logic;
signal \N__7140\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7136\ : std_logic;
signal \N__7133\ : std_logic;
signal \N__7132\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7126\ : std_logic;
signal \N__7123\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7117\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7096\ : std_logic;
signal \N__7093\ : std_logic;
signal \N__7090\ : std_logic;
signal \N__7087\ : std_logic;
signal \N__7084\ : std_logic;
signal \N__7081\ : std_logic;
signal \N__7078\ : std_logic;
signal \N__7075\ : std_logic;
signal \N__7072\ : std_logic;
signal \N__7069\ : std_logic;
signal \N__7066\ : std_logic;
signal \N__7063\ : std_logic;
signal \N__7060\ : std_logic;
signal \N__7059\ : std_logic;
signal \N__7056\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7050\ : std_logic;
signal \N__7049\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7040\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7032\ : std_logic;
signal \N__7031\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7027\ : std_logic;
signal \N__7024\ : std_logic;
signal \N__7021\ : std_logic;
signal \N__7020\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7016\ : std_logic;
signal \N__7013\ : std_logic;
signal \N__7010\ : std_logic;
signal \N__7007\ : std_logic;
signal \N__7004\ : std_logic;
signal \N__7001\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6990\ : std_logic;
signal \N__6987\ : std_logic;
signal \N__6982\ : std_logic;
signal \N__6979\ : std_logic;
signal \N__6976\ : std_logic;
signal \N__6971\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6955\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6946\ : std_logic;
signal \N__6943\ : std_logic;
signal \N__6942\ : std_logic;
signal \N__6939\ : std_logic;
signal \N__6936\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6931\ : std_logic;
signal \N__6928\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6926\ : std_logic;
signal \N__6925\ : std_logic;
signal \N__6922\ : std_logic;
signal \N__6919\ : std_logic;
signal \N__6916\ : std_logic;
signal \N__6913\ : std_logic;
signal \N__6908\ : std_logic;
signal \N__6905\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6889\ : std_logic;
signal \N__6886\ : std_logic;
signal \N__6885\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6874\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6860\ : std_logic;
signal \N__6857\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6838\ : std_logic;
signal \N__6835\ : std_logic;
signal \N__6834\ : std_logic;
signal \N__6831\ : std_logic;
signal \N__6828\ : std_logic;
signal \N__6825\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6802\ : std_logic;
signal \N__6799\ : std_logic;
signal \N__6798\ : std_logic;
signal \N__6795\ : std_logic;
signal \N__6792\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6780\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6774\ : std_logic;
signal \N__6773\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6768\ : std_logic;
signal \N__6767\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6762\ : std_logic;
signal \N__6761\ : std_logic;
signal \N__6760\ : std_logic;
signal \N__6755\ : std_logic;
signal \N__6754\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6752\ : std_logic;
signal \N__6749\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6743\ : std_logic;
signal \N__6740\ : std_logic;
signal \N__6737\ : std_logic;
signal \N__6732\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6718\ : std_logic;
signal \N__6713\ : std_logic;
signal \N__6706\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6693\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6685\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6673\ : std_logic;
signal \N__6672\ : std_logic;
signal \N__6669\ : std_logic;
signal \N__6668\ : std_logic;
signal \N__6665\ : std_logic;
signal \N__6660\ : std_logic;
signal \N__6657\ : std_logic;
signal \N__6654\ : std_logic;
signal \N__6653\ : std_logic;
signal \N__6650\ : std_logic;
signal \N__6647\ : std_logic;
signal \N__6644\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6621\ : std_logic;
signal \N__6620\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6618\ : std_logic;
signal \N__6617\ : std_logic;
signal \N__6616\ : std_logic;
signal \N__6615\ : std_logic;
signal \N__6614\ : std_logic;
signal \N__6611\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6607\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6603\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6597\ : std_logic;
signal \N__6594\ : std_logic;
signal \N__6591\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6582\ : std_logic;
signal \N__6581\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6577\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6566\ : std_logic;
signal \N__6563\ : std_logic;
signal \N__6560\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6540\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6516\ : std_logic;
signal \N__6505\ : std_logic;
signal \N__6502\ : std_logic;
signal \N__6501\ : std_logic;
signal \N__6500\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6498\ : std_logic;
signal \N__6497\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6493\ : std_logic;
signal \N__6492\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6476\ : std_logic;
signal \N__6475\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6471\ : std_logic;
signal \N__6468\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6457\ : std_logic;
signal \N__6456\ : std_logic;
signal \N__6453\ : std_logic;
signal \N__6450\ : std_logic;
signal \N__6447\ : std_logic;
signal \N__6442\ : std_logic;
signal \N__6439\ : std_logic;
signal \N__6436\ : std_logic;
signal \N__6433\ : std_logic;
signal \N__6428\ : std_logic;
signal \N__6425\ : std_logic;
signal \N__6406\ : std_logic;
signal \N__6403\ : std_logic;
signal \N__6402\ : std_logic;
signal \N__6399\ : std_logic;
signal \N__6396\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6388\ : std_logic;
signal \N__6385\ : std_logic;
signal \N__6380\ : std_logic;
signal \N__6377\ : std_logic;
signal \N__6374\ : std_logic;
signal \N__6367\ : std_logic;
signal \N__6364\ : std_logic;
signal \N__6363\ : std_logic;
signal \N__6360\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6356\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6349\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6341\ : std_logic;
signal \N__6338\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6330\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6320\ : std_logic;
signal \N__6317\ : std_logic;
signal \N__6316\ : std_logic;
signal \N__6313\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6307\ : std_logic;
signal \N__6304\ : std_logic;
signal \N__6301\ : std_logic;
signal \N__6298\ : std_logic;
signal \N__6295\ : std_logic;
signal \N__6292\ : std_logic;
signal \N__6289\ : std_logic;
signal \N__6286\ : std_logic;
signal \N__6281\ : std_logic;
signal \N__6274\ : std_logic;
signal \N__6273\ : std_logic;
signal \N__6272\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6266\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6253\ : std_logic;
signal \N__6250\ : std_logic;
signal \N__6247\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6239\ : std_logic;
signal \N__6236\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6228\ : std_logic;
signal \N__6225\ : std_logic;
signal \N__6222\ : std_logic;
signal \N__6219\ : std_logic;
signal \N__6216\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6210\ : std_logic;
signal \N__6207\ : std_logic;
signal \N__6204\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6196\ : std_logic;
signal \N__6195\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6188\ : std_logic;
signal \N__6185\ : std_logic;
signal \N__6178\ : std_logic;
signal \N__6177\ : std_logic;
signal \N__6174\ : std_logic;
signal \N__6171\ : std_logic;
signal \N__6170\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6150\ : std_logic;
signal \N__6145\ : std_logic;
signal \N__6142\ : std_logic;
signal \N__6141\ : std_logic;
signal \N__6138\ : std_logic;
signal \N__6135\ : std_logic;
signal \N__6132\ : std_logic;
signal \N__6129\ : std_logic;
signal \N__6128\ : std_logic;
signal \N__6123\ : std_logic;
signal \N__6120\ : std_logic;
signal \N__6115\ : std_logic;
signal \N__6114\ : std_logic;
signal \N__6111\ : std_logic;
signal \N__6108\ : std_logic;
signal \N__6105\ : std_logic;
signal \N__6102\ : std_logic;
signal \N__6101\ : std_logic;
signal \N__6100\ : std_logic;
signal \N__6097\ : std_logic;
signal \N__6094\ : std_logic;
signal \N__6091\ : std_logic;
signal \N__6088\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6078\ : std_logic;
signal \N__6075\ : std_logic;
signal \N__6074\ : std_logic;
signal \N__6071\ : std_logic;
signal \N__6070\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6058\ : std_logic;
signal \N__6053\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6047\ : std_logic;
signal \N__6044\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6031\ : std_logic;
signal \N__6030\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6022\ : std_logic;
signal \N__6019\ : std_logic;
signal \N__6016\ : std_logic;
signal \N__6013\ : std_logic;
signal \N__6010\ : std_logic;
signal \N__6007\ : std_logic;
signal \N__6004\ : std_logic;
signal \N__6001\ : std_logic;
signal \N__5994\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5988\ : std_logic;
signal \N__5983\ : std_logic;
signal \N__5980\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5966\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5953\ : std_logic;
signal \N__5950\ : std_logic;
signal \N__5949\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5946\ : std_logic;
signal \N__5943\ : std_logic;
signal \N__5940\ : std_logic;
signal \N__5933\ : std_logic;
signal \N__5930\ : std_logic;
signal \N__5925\ : std_logic;
signal \N__5920\ : std_logic;
signal \N__5917\ : std_logic;
signal \N__5914\ : std_logic;
signal \N__5913\ : std_logic;
signal \N__5910\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5905\ : std_logic;
signal \N__5902\ : std_logic;
signal \N__5899\ : std_logic;
signal \N__5896\ : std_logic;
signal \N__5893\ : std_logic;
signal \N__5884\ : std_logic;
signal \N__5883\ : std_logic;
signal \N__5880\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5878\ : std_logic;
signal \N__5877\ : std_logic;
signal \N__5874\ : std_logic;
signal \N__5871\ : std_logic;
signal \N__5864\ : std_logic;
signal \N__5861\ : std_logic;
signal \N__5856\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5848\ : std_logic;
signal \N__5845\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5841\ : std_logic;
signal \N__5838\ : std_logic;
signal \N__5837\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5833\ : std_logic;
signal \N__5830\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5816\ : std_logic;
signal \N__5813\ : std_logic;
signal \N__5810\ : std_logic;
signal \N__5807\ : std_logic;
signal \N__5802\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5793\ : std_logic;
signal \N__5792\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5786\ : std_logic;
signal \N__5783\ : std_logic;
signal \N__5780\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5751\ : std_logic;
signal \N__5750\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5745\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5739\ : std_logic;
signal \N__5736\ : std_logic;
signal \N__5733\ : std_logic;
signal \N__5730\ : std_logic;
signal \N__5725\ : std_logic;
signal \N__5720\ : std_logic;
signal \N__5713\ : std_logic;
signal \N__5710\ : std_logic;
signal \N__5709\ : std_logic;
signal \N__5706\ : std_logic;
signal \N__5703\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5701\ : std_logic;
signal \N__5700\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5687\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5677\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5671\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5658\ : std_logic;
signal \N__5657\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5655\ : std_logic;
signal \N__5654\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5652\ : std_logic;
signal \N__5651\ : std_logic;
signal \N__5650\ : std_logic;
signal \N__5649\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5647\ : std_logic;
signal \N__5646\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5642\ : std_logic;
signal \N__5641\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5639\ : std_logic;
signal \N__5638\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5636\ : std_logic;
signal \N__5635\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5633\ : std_logic;
signal \N__5632\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5630\ : std_logic;
signal \N__5629\ : std_logic;
signal \N__5628\ : std_logic;
signal \N__5627\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5625\ : std_logic;
signal \N__5624\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5533\ : std_logic;
signal \N__5530\ : std_logic;
signal \N__5527\ : std_logic;
signal \N__5524\ : std_logic;
signal \N__5521\ : std_logic;
signal \N__5520\ : std_logic;
signal \N__5517\ : std_logic;
signal \N__5516\ : std_logic;
signal \N__5513\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5502\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5485\ : std_logic;
signal \N__5484\ : std_logic;
signal \N__5481\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5467\ : std_logic;
signal \N__5464\ : std_logic;
signal \N__5461\ : std_logic;
signal \N__5458\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5451\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5442\ : std_logic;
signal \N__5439\ : std_logic;
signal \N__5436\ : std_logic;
signal \N__5433\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5421\ : std_logic;
signal \N__5420\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5418\ : std_logic;
signal \N__5417\ : std_logic;
signal \N__5416\ : std_logic;
signal \N__5415\ : std_logic;
signal \N__5414\ : std_logic;
signal \N__5413\ : std_logic;
signal \N__5410\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5395\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5376\ : std_logic;
signal \N__5373\ : std_logic;
signal \N__5370\ : std_logic;
signal \N__5367\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5358\ : std_logic;
signal \N__5357\ : std_logic;
signal \N__5356\ : std_logic;
signal \N__5353\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5349\ : std_logic;
signal \N__5346\ : std_logic;
signal \N__5343\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5341\ : std_logic;
signal \N__5340\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5336\ : std_logic;
signal \N__5331\ : std_logic;
signal \N__5328\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5315\ : std_logic;
signal \N__5302\ : std_logic;
signal \N__5301\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5298\ : std_logic;
signal \N__5297\ : std_logic;
signal \N__5294\ : std_logic;
signal \N__5289\ : std_logic;
signal \N__5284\ : std_logic;
signal \N__5283\ : std_logic;
signal \N__5280\ : std_logic;
signal \N__5277\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5269\ : std_logic;
signal \N__5266\ : std_logic;
signal \N__5261\ : std_logic;
signal \N__5258\ : std_logic;
signal \N__5255\ : std_logic;
signal \N__5250\ : std_logic;
signal \N__5245\ : std_logic;
signal \N__5244\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5242\ : std_logic;
signal \N__5241\ : std_logic;
signal \N__5238\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5226\ : std_logic;
signal \N__5221\ : std_logic;
signal \N__5214\ : std_logic;
signal \N__5209\ : std_logic;
signal \N__5206\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5200\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5194\ : std_logic;
signal \N__5193\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5186\ : std_logic;
signal \N__5183\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5181\ : std_logic;
signal \N__5178\ : std_logic;
signal \N__5175\ : std_logic;
signal \N__5172\ : std_logic;
signal \N__5171\ : std_logic;
signal \N__5168\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5160\ : std_logic;
signal \N__5157\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5149\ : std_logic;
signal \N__5146\ : std_logic;
signal \N__5143\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5131\ : std_logic;
signal \N__5128\ : std_logic;
signal \N__5125\ : std_logic;
signal \N__5124\ : std_logic;
signal \N__5121\ : std_logic;
signal \N__5118\ : std_logic;
signal \N__5113\ : std_logic;
signal \N__5110\ : std_logic;
signal \N__5107\ : std_logic;
signal \N__5104\ : std_logic;
signal \N__5101\ : std_logic;
signal \N__5100\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5086\ : std_logic;
signal \N__5083\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5081\ : std_logic;
signal \N__5080\ : std_logic;
signal \N__5077\ : std_logic;
signal \N__5074\ : std_logic;
signal \N__5069\ : std_logic;
signal \N__5064\ : std_logic;
signal \N__5061\ : std_logic;
signal \N__5058\ : std_logic;
signal \N__5047\ : std_logic;
signal \N__5044\ : std_logic;
signal \N__5041\ : std_logic;
signal \N__5038\ : std_logic;
signal \N__5035\ : std_logic;
signal \N__5032\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5028\ : std_logic;
signal \N__5025\ : std_logic;
signal \N__5022\ : std_logic;
signal \N__5021\ : std_logic;
signal \N__5016\ : std_logic;
signal \N__5013\ : std_logic;
signal \N__5012\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__4996\ : std_logic;
signal \N__4993\ : std_logic;
signal \N__4990\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4988\ : std_logic;
signal \N__4983\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4979\ : std_logic;
signal \N__4978\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4974\ : std_logic;
signal \N__4971\ : std_logic;
signal \N__4968\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4962\ : std_logic;
signal \N__4959\ : std_logic;
signal \N__4954\ : std_logic;
signal \N__4951\ : std_logic;
signal \N__4936\ : std_logic;
signal \N__4933\ : std_logic;
signal \N__4932\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4930\ : std_logic;
signal \N__4929\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4917\ : std_logic;
signal \N__4914\ : std_logic;
signal \N__4911\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4909\ : std_logic;
signal \N__4908\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4906\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4893\ : std_logic;
signal \N__4888\ : std_logic;
signal \N__4881\ : std_logic;
signal \N__4870\ : std_logic;
signal \N__4869\ : std_logic;
signal \N__4866\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4864\ : std_logic;
signal \N__4863\ : std_logic;
signal \N__4860\ : std_logic;
signal \N__4857\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4843\ : std_logic;
signal \N__4842\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4840\ : std_logic;
signal \N__4839\ : std_logic;
signal \N__4836\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4830\ : std_logic;
signal \N__4827\ : std_logic;
signal \N__4824\ : std_logic;
signal \N__4813\ : std_logic;
signal \N__4810\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4771\ : std_logic;
signal \N__4768\ : std_logic;
signal \N__4767\ : std_logic;
signal \N__4764\ : std_logic;
signal \N__4761\ : std_logic;
signal \N__4760\ : std_logic;
signal \N__4759\ : std_logic;
signal \N__4758\ : std_logic;
signal \N__4757\ : std_logic;
signal \N__4754\ : std_logic;
signal \N__4751\ : std_logic;
signal \N__4746\ : std_logic;
signal \N__4743\ : std_logic;
signal \N__4740\ : std_logic;
signal \N__4739\ : std_logic;
signal \N__4738\ : std_logic;
signal \N__4737\ : std_logic;
signal \N__4736\ : std_logic;
signal \N__4733\ : std_logic;
signal \N__4730\ : std_logic;
signal \N__4727\ : std_logic;
signal \N__4714\ : std_logic;
signal \N__4705\ : std_logic;
signal \N__4704\ : std_logic;
signal \N__4703\ : std_logic;
signal \N__4702\ : std_logic;
signal \N__4701\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4689\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4685\ : std_logic;
signal \N__4684\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4677\ : std_logic;
signal \N__4674\ : std_logic;
signal \N__4671\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4642\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4638\ : std_logic;
signal \N__4635\ : std_logic;
signal \N__4630\ : std_logic;
signal \N__4627\ : std_logic;
signal \N__4624\ : std_logic;
signal \N__4621\ : std_logic;
signal \N__4618\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4612\ : std_logic;
signal \N__4609\ : std_logic;
signal \N__4606\ : std_logic;
signal \N__4603\ : std_logic;
signal \N__4600\ : std_logic;
signal \N__4597\ : std_logic;
signal \N__4594\ : std_logic;
signal \N__4591\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4585\ : std_logic;
signal \N__4582\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4575\ : std_logic;
signal \N__4572\ : std_logic;
signal \N__4569\ : std_logic;
signal \N__4564\ : std_logic;
signal \N__4561\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4554\ : std_logic;
signal \N__4551\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4545\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4537\ : std_logic;
signal \N__4534\ : std_logic;
signal \N__4531\ : std_logic;
signal \N__4528\ : std_logic;
signal \N__4525\ : std_logic;
signal \N__4524\ : std_logic;
signal \N__4521\ : std_logic;
signal \N__4518\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4510\ : std_logic;
signal \N__4507\ : std_logic;
signal \N__4504\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4500\ : std_logic;
signal \N__4499\ : std_logic;
signal \N__4496\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4490\ : std_logic;
signal \N__4487\ : std_logic;
signal \N__4480\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4478\ : std_logic;
signal \N__4475\ : std_logic;
signal \N__4472\ : std_logic;
signal \N__4469\ : std_logic;
signal \N__4468\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4466\ : std_logic;
signal \N__4463\ : std_logic;
signal \N__4460\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4451\ : std_logic;
signal \N__4448\ : std_logic;
signal \N__4443\ : std_logic;
signal \N__4438\ : std_logic;
signal \N__4435\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4423\ : std_logic;
signal \N__4420\ : std_logic;
signal \N__4419\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4416\ : std_logic;
signal \N__4415\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4409\ : std_logic;
signal \N__4406\ : std_logic;
signal \N__4401\ : std_logic;
signal \N__4400\ : std_logic;
signal \N__4399\ : std_logic;
signal \N__4398\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4396\ : std_logic;
signal \N__4393\ : std_logic;
signal \N__4390\ : std_logic;
signal \N__4385\ : std_logic;
signal \N__4382\ : std_logic;
signal \N__4371\ : std_logic;
signal \N__4368\ : std_logic;
signal \N__4357\ : std_logic;
signal \N__4354\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4342\ : std_logic;
signal \N__4341\ : std_logic;
signal \N__4338\ : std_logic;
signal \N__4335\ : std_logic;
signal \N__4330\ : std_logic;
signal \N__4327\ : std_logic;
signal \N__4326\ : std_logic;
signal \N__4321\ : std_logic;
signal \N__4320\ : std_logic;
signal \N__4317\ : std_logic;
signal \N__4314\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4306\ : std_logic;
signal \N__4303\ : std_logic;
signal \N__4300\ : std_logic;
signal \N__4297\ : std_logic;
signal \N__4296\ : std_logic;
signal \N__4293\ : std_logic;
signal \N__4290\ : std_logic;
signal \N__4285\ : std_logic;
signal \N__4282\ : std_logic;
signal \N__4279\ : std_logic;
signal \N__4276\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4270\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4261\ : std_logic;
signal \N__4258\ : std_logic;
signal \N__4255\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4246\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4240\ : std_logic;
signal \N__4239\ : std_logic;
signal \N__4236\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4224\ : std_logic;
signal \N__4223\ : std_logic;
signal \N__4220\ : std_logic;
signal \N__4215\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4201\ : std_logic;
signal \N__4200\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4177\ : std_logic;
signal \N__4174\ : std_logic;
signal \N__4171\ : std_logic;
signal \N__4168\ : std_logic;
signal \N__4165\ : std_logic;
signal \N__4162\ : std_logic;
signal \N__4159\ : std_logic;
signal \N__4156\ : std_logic;
signal \N__4153\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4144\ : std_logic;
signal \N__4143\ : std_logic;
signal \N__4142\ : std_logic;
signal \N__4139\ : std_logic;
signal \N__4138\ : std_logic;
signal \N__4137\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4128\ : std_logic;
signal \N__4127\ : std_logic;
signal \N__4124\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4116\ : std_logic;
signal \N__4113\ : std_logic;
signal \N__4110\ : std_logic;
signal \N__4107\ : std_logic;
signal \N__4104\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4102\ : std_logic;
signal \N__4101\ : std_logic;
signal \N__4098\ : std_logic;
signal \N__4095\ : std_logic;
signal \N__4092\ : std_logic;
signal \N__4087\ : std_logic;
signal \N__4080\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4062\ : std_logic;
signal \N__4045\ : std_logic;
signal \N__4044\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4042\ : std_logic;
signal \N__4039\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4024\ : std_logic;
signal \N__4023\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4021\ : std_logic;
signal \N__4020\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4014\ : std_logic;
signal \N__4011\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__3996\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3978\ : std_logic;
signal \N__3975\ : std_logic;
signal \N__3972\ : std_logic;
signal \N__3969\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3961\ : std_logic;
signal \N__3958\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3934\ : std_logic;
signal \N__3931\ : std_logic;
signal \N__3928\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3924\ : std_logic;
signal \N__3923\ : std_logic;
signal \N__3920\ : std_logic;
signal \N__3915\ : std_logic;
signal \N__3910\ : std_logic;
signal \N__3907\ : std_logic;
signal \N__3904\ : std_logic;
signal \N__3901\ : std_logic;
signal \N__3898\ : std_logic;
signal \N__3895\ : std_logic;
signal \N__3892\ : std_logic;
signal \N__3891\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3884\ : std_logic;
signal \N__3883\ : std_logic;
signal \N__3880\ : std_logic;
signal \N__3877\ : std_logic;
signal \N__3874\ : std_logic;
signal \N__3871\ : std_logic;
signal \N__3868\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3856\ : std_logic;
signal \N__3855\ : std_logic;
signal \N__3850\ : std_logic;
signal \N__3849\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3847\ : std_logic;
signal \N__3844\ : std_logic;
signal \N__3841\ : std_logic;
signal \N__3838\ : std_logic;
signal \N__3835\ : std_logic;
signal \N__3826\ : std_logic;
signal \N__3823\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3811\ : std_logic;
signal \N__3810\ : std_logic;
signal \N__3807\ : std_logic;
signal \N__3804\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3798\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3778\ : std_logic;
signal \N__3777\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3771\ : std_logic;
signal \N__3768\ : std_logic;
signal \N__3765\ : std_logic;
signal \N__3760\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3754\ : std_logic;
signal \N__3751\ : std_logic;
signal \N__3748\ : std_logic;
signal \N__3745\ : std_logic;
signal \N__3742\ : std_logic;
signal \N__3739\ : std_logic;
signal \N__3736\ : std_logic;
signal \N__3733\ : std_logic;
signal \N__3732\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3716\ : std_logic;
signal \N__3709\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3703\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3697\ : std_logic;
signal \N__3694\ : std_logic;
signal \N__3691\ : std_logic;
signal \N__3688\ : std_logic;
signal \N__3685\ : std_logic;
signal \N__3682\ : std_logic;
signal \N__3679\ : std_logic;
signal \N__3676\ : std_logic;
signal \N__3673\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3664\ : std_logic;
signal \N__3661\ : std_logic;
signal \N__3658\ : std_logic;
signal \N__3655\ : std_logic;
signal \N__3652\ : std_logic;
signal \N__3649\ : std_logic;
signal \N__3648\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3642\ : std_logic;
signal \N__3639\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3628\ : std_logic;
signal \N__3627\ : std_logic;
signal \N__3624\ : std_logic;
signal \N__3621\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3613\ : std_logic;
signal \N__3610\ : std_logic;
signal \N__3607\ : std_logic;
signal \N__3604\ : std_logic;
signal \N__3601\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3595\ : std_logic;
signal \N__3592\ : std_logic;
signal \N__3589\ : std_logic;
signal \N__3588\ : std_logic;
signal \N__3585\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3573\ : std_logic;
signal \N__3570\ : std_logic;
signal \N__3565\ : std_logic;
signal \N__3562\ : std_logic;
signal \N__3559\ : std_logic;
signal \N__3558\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3553\ : std_logic;
signal \N__3552\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3548\ : std_logic;
signal \N__3545\ : std_logic;
signal \N__3544\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3531\ : std_logic;
signal \N__3528\ : std_logic;
signal \N__3525\ : std_logic;
signal \N__3522\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3512\ : std_logic;
signal \N__3507\ : std_logic;
signal \N__3502\ : std_logic;
signal \N__3499\ : std_logic;
signal \N__3496\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3490\ : std_logic;
signal \N__3487\ : std_logic;
signal \N__3484\ : std_logic;
signal \N__3481\ : std_logic;
signal \N__3478\ : std_logic;
signal \N__3475\ : std_logic;
signal \N__3472\ : std_logic;
signal \N__3469\ : std_logic;
signal \N__3466\ : std_logic;
signal \N__3463\ : std_logic;
signal \N__3460\ : std_logic;
signal \N__3457\ : std_logic;
signal \N__3454\ : std_logic;
signal \N__3451\ : std_logic;
signal \N__3448\ : std_logic;
signal \N__3445\ : std_logic;
signal \N__3444\ : std_logic;
signal \N__3439\ : std_logic;
signal \N__3436\ : std_logic;
signal \N__3433\ : std_logic;
signal \N__3430\ : std_logic;
signal \N__3427\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3415\ : std_logic;
signal \N__3412\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3403\ : std_logic;
signal \N__3400\ : std_logic;
signal \N__3397\ : std_logic;
signal \N__3394\ : std_logic;
signal \N__3391\ : std_logic;
signal \N__3388\ : std_logic;
signal \N__3385\ : std_logic;
signal \N__3382\ : std_logic;
signal \N__3379\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3373\ : std_logic;
signal \N__3370\ : std_logic;
signal \N__3367\ : std_logic;
signal \N__3364\ : std_logic;
signal \N__3361\ : std_logic;
signal \N__3358\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3349\ : std_logic;
signal \N__3346\ : std_logic;
signal \N__3343\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3337\ : std_logic;
signal \N__3334\ : std_logic;
signal \N__3331\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3325\ : std_logic;
signal \N__3322\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3318\ : std_logic;
signal \N__3315\ : std_logic;
signal \N__3312\ : std_logic;
signal \N__3309\ : std_logic;
signal \N__3306\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3288\ : std_logic;
signal \N__3285\ : std_logic;
signal \N__3282\ : std_logic;
signal \N__3277\ : std_logic;
signal \N__3274\ : std_logic;
signal \N__3271\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3265\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3259\ : std_logic;
signal \N__3256\ : std_logic;
signal \N__3253\ : std_logic;
signal \N__3250\ : std_logic;
signal \N__3247\ : std_logic;
signal \N__3244\ : std_logic;
signal \N__3241\ : std_logic;
signal \N__3238\ : std_logic;
signal \N__3235\ : std_logic;
signal \N__3232\ : std_logic;
signal \N__3229\ : std_logic;
signal \N__3226\ : std_logic;
signal \VCCG0\ : std_logic;
signal \GNDG0\ : std_logic;
signal \G_138\ : std_logic;
signal \G_138_cascade_\ : std_logic;
signal \uut.buf_clk_1\ : std_logic;
signal \INVuut.b_reg.ff6.qC_net\ : std_logic;
signal \INVuut.b_reg.ff7.qC_net\ : std_logic;
signal \INVuut.acc.ff2.qC_net\ : std_logic;
signal \uut.AR_BUF.out_1_1_iv_3_1Z0Z_0_cascade_\ : std_logic;
signal \uut.AR_BUF.out_1_1_ivZ0Z_0_cascade_\ : std_logic;
signal \uut.out_1_1_iv_2_cascade_\ : std_logic;
signal \INVuut.AR.ff2.qC_net\ : std_logic;
signal \uut.ALU_main.N_47_cascade_\ : std_logic;
signal \uut.seq.un1_HLT_1_reti_cascade_\ : std_logic;
signal \uut.un1_HLT_0\ : std_logic;
signal \INVuut.seq.q_ret_1C_net\ : std_logic;
signal \uut.ALU_main.N_46_cascade_\ : std_logic;
signal \uut.alu_out_m_5_cascade_\ : std_logic;
signal \uut.bus_5_cascade_\ : std_logic;
signal \uut.alu_out_m_7_cascade_\ : std_logic;
signal \INVuut.b_reg.ff8.qC_net\ : std_logic;
signal \uut.acc_out_m_7_cascade_\ : std_logic;
signal \uut.bus_7_cascade_\ : std_logic;
signal \uut.N_1_0\ : std_logic;
signal \LED5_c\ : std_logic;
signal \INVuut.out_reg.ff5.qC_net\ : std_logic;
signal \uut.out_1_2_iv_3_cascade_\ : std_logic;
signal \LED1_c\ : std_logic;
signal \INVuut.out_reg.ff1.qC_net\ : std_logic;
signal \INVuut.acc.ff3.qC_net\ : std_logic;
signal \uut.program_counter_m_2_cascade_\ : std_logic;
signal \uut.AR_BUF.N_8\ : std_logic;
signal \uut.program_counter_m_2\ : std_logic;
signal \uut.AR_BUF.g0_0_0Z0Z_1\ : std_logic;
signal \uut.out_1_0_ivdup_2_cascade_\ : std_logic;
signal \uut.ALU_main.N_43\ : std_logic;
signal \uut.ir_out_m_d_1\ : std_logic;
signal \uut.bus_6_cascade_\ : std_logic;
signal \uut.q_RNIDGA71_cascade_\ : std_logic;
signal \INVuut.b_reg.ff5.qC_net\ : std_logic;
signal \uut.ALU_main.N_45_cascade_\ : std_logic;
signal \uut.alu_out_m_4_cascade_\ : std_logic;
signal \uut.data_1_2_ivdup_cascade_\ : std_logic;
signal \uut.N_4_0\ : std_logic;
signal \uut.data_1_2_iv_0\ : std_logic;
signal \uut.b_reg_out_4\ : std_logic;
signal \INVuut.IR.ff5.q_0_neC_net\ : std_logic;
signal \uut.AR_BUF.out_1_0_iv_2Z0Z_0\ : std_logic;
signal \uut.ir_out_m_d_2_cascade_\ : std_logic;
signal \INVuut.seq.q_retC_net\ : std_logic;
signal \uut.ALU_main.N_48\ : std_logic;
signal \uut.AR_BUF.out_1_0_iv_2_1Z0Z_1\ : std_logic;
signal \INVuut.IR.ff1.q_neC_net\ : std_logic;
signal \uut.AR_BUF.g0_0_a5_0Z0Z_2_cascade_\ : std_logic;
signal \uut.AR_BUF.N_9\ : std_logic;
signal \uut.AR_BUF.g0_1_a10_3Z0Z_2\ : std_logic;
signal \uut.AR_BUF.g0_0_o5_0Z0Z_0\ : std_logic;
signal \uut.AR_BUF.g0_1_a10_3_cascade_\ : std_logic;
signal \uut.AR_BUF.N_7\ : std_logic;
signal \uut.AR_BUF.N_13_cascade_\ : std_logic;
signal \uut.AR_BUF.g0_1_0Z0Z_5_cascade_\ : std_logic;
signal \uut.AR_BUF.g0_1_0Z0Z_1\ : std_logic;
signal \uut.AR_out_1\ : std_logic;
signal \uut.AR_BUF.g0_1_0_4_0\ : std_logic;
signal \uut.ir_out_1\ : std_logic;
signal \uut.AR_BUF.N_10\ : std_logic;
signal \uut.AR_BUF.g0_1_0_0_0\ : std_logic;
signal \uut.ir_out_m_d_0\ : std_logic;
signal \uut.pc.N_4_i_1_cascade_\ : std_logic;
signal \uut.alu_out_m_2\ : std_logic;
signal \INVuut.b_reg.ff3.qC_net\ : std_logic;
signal \uut.ALU_main.N_43_0_cascade_\ : std_logic;
signal \uut.T_1_fast_RNIVM0N3_0_cascade_\ : std_logic;
signal \uut.pc.N_11\ : std_logic;
signal \uut.seq.counter.T_2_rep1_RNI8TEZ0Z81_cascade_\ : std_logic;
signal \uut.seq.counter.un2_MAR_LD_cascade_\ : std_logic;
signal \uut.D_1_0_cascade_\ : std_logic;
signal \uut.seq.q_ret_RNI52E81Z0Z_0\ : std_logic;
signal \uut.T_2_rep1_RNI6BLF1_cascade_\ : std_logic;
signal \uut.un17_IR_OE_0\ : std_logic;
signal \uut.IR.ir_out_m_c_d_1_3_cascade_\ : std_logic;
signal \uut.ir_out_m_c_d_3_cascade_\ : std_logic;
signal \INVuut.IR.ff4.q_neC_net\ : std_logic;
signal \uut.seq.counter.T_2_rep1_RNIGC8CZ0Z1\ : std_logic;
signal \uut.seq.un13_ACC_LD_xZ0Z1_cascade_\ : std_logic;
signal \uut.un1_HLT_1\ : std_logic;
signal \uut.N_5_0\ : std_logic;
signal \uut.bus_6\ : std_logic;
signal \INVuut.IR.ff7.q_ret_1_fastC_net\ : std_logic;
signal \uut.bus_7\ : std_logic;
signal \uut.seq.D_2_0_x_cascade_\ : std_logic;
signal \uut.q_0_fast\ : std_logic;
signal \uut.data_1_2_ivdup\ : std_logic;
signal \INVuut.IR.ff5.q_0_rep1C_net\ : std_logic;
signal \uut.seq.counter.un4_ACC_LD_cascade_\ : std_logic;
signal \uut.seq.counter.ACC_LD_0_0\ : std_logic;
signal \uut.N_2_0\ : std_logic;
signal \INVuut.seq.counter.T_1_fast_3C_net\ : std_logic;
signal \uut.q_ret_1_fast_0\ : std_logic;
signal \uut.AR_BUF.g0_3Z0Z_3_cascade_\ : std_logic;
signal \INVuut.acc.ff1.qC_net\ : std_logic;
signal \uut.AR_BUF.out_1_2_ivZ0Z_1\ : std_logic;
signal \uut.ir_out_7\ : std_logic;
signal \uut.ir_out_6\ : std_logic;
signal \uut.AR_BUF.g0_3_a10_1Z0Z_1\ : std_logic;
signal \uut.D_1_0\ : std_logic;
signal \uut.AR_BUF.g0_3_a10_0Z0Z_2_cascade_\ : std_logic;
signal \uut.AR_BUF.g0_3Z0Z_0\ : std_logic;
signal \uut.ir_out_m_c_d_0_cascade_\ : std_logic;
signal \uut.AR_BUF.out_1_2_ivZ0Z_2\ : std_logic;
signal \uut.AR_BUF.g0_1_a10_4Z0Z_1\ : std_logic;
signal \uut.AR_BUF.g0_3Z0Z_2_cascade_\ : std_logic;
signal \uut.AR_BUF.g0_3Z0Z_6_cascade_\ : std_logic;
signal \INVuut.AR.ff1.q_neC_net\ : std_logic;
signal \uut.AR_out_0\ : std_logic;
signal \uut.T_1_RNIVVKI3_3\ : std_logic;
signal \uut.program_counter_m_0\ : std_logic;
signal \uut.pc.G_26_i_a4_5_sx_cascade_\ : std_logic;
signal \uut.pc.G_26_i_a4_5\ : std_logic;
signal \uut.ir_out_m_c_c_0\ : std_logic;
signal \uut.alu_out_m_0_0\ : std_logic;
signal \uut.alu_out_m_0\ : std_logic;
signal \INVuut.b_reg.ff4.qC_net\ : std_logic;
signal \uut.pc.program_counter_4_a1_0_0_1_cascade_\ : std_logic;
signal \uut.pc.g2_0\ : std_logic;
signal \uut.pc.N_77_0\ : std_logic;
signal \uut.pc.g1_0_cascade_\ : std_logic;
signal \uut.pc.program_counter_0_1_1\ : std_logic;
signal \uut.S0_0_i\ : std_logic;
signal \bfn_9_12_0_\ : std_logic;
signal \uut.un1_A_cry_0_s\ : std_logic;
signal \uut.ALU_main.un1_A_cry_0_c_THRU_CO\ : std_logic;
signal \uut.ALU_main.un1_A_cry_0\ : std_logic;
signal \uut.ALU_main.un1_A_cry_1_c_RNI7KLZ0Z45\ : std_logic;
signal \uut.ALU_main.un1_A_cry_1\ : std_logic;
signal \uut.ALU_main.un1_A_axb_3_l_ofxZ0\ : std_logic;
signal \uut.ALU_main.un1_A_cry_2_cZ0\ : std_logic;
signal \uut.ALU_main.un1_A_axb_4_l_ofxZ0\ : std_logic;
signal \uut.ALU_main.un1_A_cry_3_c_RNIF4UZ0Z45\ : std_logic;
signal \uut.ALU_main.un1_A_cry_3\ : std_logic;
signal \uut.ALU_main.un1_A_cry_4_c_RNIJCZ0Z255\ : std_logic;
signal \uut.ALU_main.un1_A_cry_4\ : std_logic;
signal \uut.ALU_main.un1_A_cry_5_c_RNINKZ0Z655\ : std_logic;
signal \uut.ALU_main.un1_A_cry_5\ : std_logic;
signal \uut.ALU_main.un1_A_cry_6\ : std_logic;
signal \bfn_9_13_0_\ : std_logic;
signal \uut.ALU_main.un1_A_cry_6_c_RNINIMNZ0Z4\ : std_logic;
signal \uut.ALU_main.un1_A_axb_1_l_ofxZ0\ : std_logic;
signal \uut.b_reg_out_6\ : std_logic;
signal \uut.ALU_main.un1_A_axb_6_l_ofxZ0\ : std_logic;
signal \uut.b_reg_out_5\ : std_logic;
signal \uut.ALU_main.un1_A_axb_5_l_ofxZ0\ : std_logic;
signal \uut.ALU_main.un1_A_axb_0_l_ofxZ0\ : std_logic;
signal \uut.b_reg_out_7\ : std_logic;
signal \uut.ALU_main.un1_A_axbZ0Z_7\ : std_logic;
signal \uut.b_reg_out_2\ : std_logic;
signal \uut.acc_out_2\ : std_logic;
signal \uut.un13_ACC_LD\ : std_logic;
signal \uut.ALU_main.un1_A_axb_2_l_ofxZ0\ : std_logic;
signal \uut.seq.counter.T_2_rep1_RNIJDGJZ0_cascade_\ : std_logic;
signal \uut.seq.D_4\ : std_logic;
signal \uut.D_1_3_cascade_\ : std_logic;
signal \uut.un7_ACC_LD\ : std_logic;
signal \uut.ir_out_4\ : std_logic;
signal \uut.seq.counter.T_1_fastZ0Z_3\ : std_logic;
signal \uut.seq.counter.T_4_cascade_\ : std_logic;
signal \uut.seq.counter.T_1_fast_RNI4JTR1_0Z0Z_0\ : std_logic;
signal \uut.T_2_rep1\ : std_logic;
signal \uut.seq.counter.T_2_rep1_RNIV9NUZ0\ : std_logic;
signal \uut.bus_5\ : std_logic;
signal \uut.q_0_fast_1\ : std_logic;
signal \uut.seq.counter.T_1_fastZ0Z_0\ : std_logic;
signal \INVuut.IR.ff6.q_0_fastC_net\ : std_logic;
signal \uut.ir_out_fast_4\ : std_logic;
signal \uut.ir_out_5\ : std_logic;
signal \uut.q_ret_1_fast\ : std_logic;
signal \uut.seq.counter.T_4\ : std_logic;
signal \uut.seq.un10_ACC_LD_xZ0Z1_cascade_\ : std_logic;
signal \uut.T_1_fast_RNI28LI1_0_cascade_\ : std_logic;
signal \uut.N_41\ : std_logic;
signal \uut.q_0_fast_0\ : std_logic;
signal \uut.seq.counter.T_fastZ0Z_2\ : std_logic;
signal \uut.seq.counter.T_fast_RNIH09PZ0Z_2_cascade_\ : std_logic;
signal \uut.ir_out_4_rep1\ : std_logic;
signal \uut.ir_out_0\ : std_logic;
signal \uut.acc_out_0\ : std_logic;
signal \uut.OUT_LD_cascade_\ : std_logic;
signal \uut.pc.G_26_i_a4_1\ : std_logic;
signal \uut.acc_out_1\ : std_logic;
signal \uut.ALU_main.ALU_Out_0Z0Z_1_cascade_\ : std_logic;
signal \uut.un1_A_cry_0_c_RNI3CH45\ : std_logic;
signal \INVuut.seq.counter.T_1_4C_net\ : std_logic;
signal \uut.seq.counter.un2_MAR_LD\ : std_logic;
signal \uut.pc.g1\ : std_logic;
signal \uut.pc.un1_inc_0_0_cascade_\ : std_logic;
signal \INVuut.seq.counter.T_1_1C_net\ : std_logic;
signal \uut.un17_IR_OE\ : std_logic;
signal \uut.PC_LD_0_0\ : std_logic;
signal \uut.PC_LD_0_0_cascade_\ : std_logic;
signal \uut.pc.un1_inc_0\ : std_logic;
signal \uut.pc.un1_inc_0_cascade_\ : std_logic;
signal \uut.pc.program_counter_4_1_2\ : std_logic;
signal \uut.m13\ : std_logic;
signal \INVuut.mar.ff2.q_neC_net\ : std_logic;
signal \uut.program_counter_2\ : std_logic;
signal \uut.program_counter_1\ : std_logic;
signal \uut.program_counter_0\ : std_logic;
signal \uut.pc.program_counter_RNO_1Z0Z_2\ : std_logic;
signal \uut.N_44_0_cascade_\ : std_logic;
signal \uut.pc.g0_rn_1\ : std_logic;
signal \uut.pc.alu_out_m_0_3_cascade_\ : std_logic;
signal \uut.buf_clk_1_g\ : std_logic;
signal \uut.ALU_main.N_44_1\ : std_logic;
signal \uut.T_1_fast_RNI28LI1_0\ : std_logic;
signal \uut.b_reg_out_3\ : std_logic;
signal \uut.un1_A_cry_2_c_RNIBSP45\ : std_logic;
signal \uut.un1_ALU_en_0\ : std_logic;
signal \uut.ALU_main.N_44_cascade_\ : std_logic;
signal \uut.T_1_fast_RNIVM0N3_0\ : std_logic;
signal \uut.acc_out_m_6\ : std_logic;
signal \uut.alu_out_m_6\ : std_logic;
signal \uut.mem.N_29_mux\ : std_logic;
signal \uut.acc_out_6\ : std_logic;
signal \uut.acc_out_m_7\ : std_logic;
signal \uut.alu_out_m_7\ : std_logic;
signal \uut.acc_out_7\ : std_logic;
signal \uut.alu_out_m_5\ : std_logic;
signal \uut.acc_out_m_5\ : std_logic;
signal \uut.mem.m20\ : std_logic;
signal \uut.acc_out_5\ : std_logic;
signal \uut.q_RNIDGA71\ : std_logic;
signal \uut.mem.i2_mux\ : std_logic;
signal \uut.alu_out_m_4\ : std_logic;
signal \uut.acc_out_4\ : std_logic;
signal \INVuut.acc.ff4.qC_net\ : std_logic;
signal \uut.ACC_LD_0_i\ : std_logic;
signal \uut.seq.D_2_1\ : std_logic;
signal \uut.ir_out_i_2_6\ : std_logic;
signal \uut.seq.D_2\ : std_logic;
signal \uut.ir_out_i_2_5\ : std_logic;
signal \uut.B_LD_0_1_tz_cascade_\ : std_logic;
signal \uut.mem.i2_mux_0\ : std_logic;
signal \uut.out_1_0_iv_2_1\ : std_logic;
signal \LED3_c\ : std_logic;
signal \INVuut.out_reg.ff3.qC_net\ : std_logic;
signal \uut.m10\ : std_logic;
signal \uut.m10_cascade_\ : std_logic;
signal \uut.b_reg_out_0\ : std_logic;
signal \uut.alu_out_m_1\ : std_logic;
signal \uut.N_11_i_m\ : std_logic;
signal \uut.out_1_1_iv_3dup_1\ : std_logic;
signal \uut.b_reg_out_1\ : std_logic;
signal \INVuut.b_reg.ff1.qC_net\ : std_logic;
signal \uut.B_LD_0_i\ : std_logic;
signal \uut.inc\ : std_logic;
signal \uut.ir_out_2\ : std_logic;
signal \INVuut.IR.ff3.qC_net\ : std_logic;
signal \uut.N_14_0\ : std_logic;
signal \uut.alu_out_m_0_2\ : std_logic;
signal \uut.out_1_0_iv_3_cascade_\ : std_logic;
signal \uut.AR_out_2\ : std_logic;
signal \INVuut.AR.ff3.qC_net\ : std_logic;
signal \uut.un11_MAR_LD\ : std_logic;
signal \uut.MAR_LD_1\ : std_logic;
signal \uut.seq.counter.MAR_LD_0_0\ : std_logic;
signal \uut.MAR_LD_1_cascade_\ : std_logic;
signal \uut.N_16_0\ : std_logic;
signal \uut.alu_out_m_1_3\ : std_logic;
signal \uut.AR_BUF.g0Z0Z_5_cascade_\ : std_logic;
signal \INVuut.AR.ff4.q_neC_net\ : std_logic;
signal \uut.AR_LD\ : std_logic;
signal \uut.un14_MAR_LD\ : std_logic;
signal \uut.un8_MAR_LD\ : std_logic;
signal \uut.un1_IR_OE_4_1\ : std_logic;
signal \uut.pc.un1_inc_0_0\ : std_logic;
signal \uut.ir_out_m_d_3_cascade_\ : std_logic;
signal \uut.pc.g0_sn\ : std_logic;
signal \uut.seq.counter.T_1Z0Z_4\ : std_logic;
signal \INVuut.seq.counter.T_1_0C_net\ : std_logic;
signal \uut.AR_BUF.out_1_ivdupZ0Z_0_cascade_\ : std_logic;
signal \uut.g0_0\ : std_logic;
signal \uut.AR_out_3\ : std_logic;
signal \uut.g1_cascade_\ : std_logic;
signal \uut.T_2_rep1_RNI6BLF1\ : std_logic;
signal \uut.AR_BUF.g0_1_0\ : std_logic;
signal \uut.T_2\ : std_logic;
signal \uut.T_0\ : std_logic;
signal \uut.program_counter_3\ : std_logic;
signal \uut.D_6\ : std_logic;
signal \uut.program_counter_m_3\ : std_logic;
signal \uut.acc_out_3\ : std_logic;
signal \uut.ir_out_3\ : std_logic;
signal \uut.un5_MAR_LD\ : std_logic;
signal \uut.AR_BUF.out_1_ivZ0Z_0_cascade_\ : std_logic;
signal \uut.out_1_iv_2\ : std_logic;
signal \uut.out_1_iv_2_1_cascade_\ : std_logic;
signal \uut.OUT_LD\ : std_logic;
signal \LED4_c\ : std_logic;
signal \uut.alu_out_m_3\ : std_logic;
signal \uut.m15_cascade_\ : std_logic;
signal \uut.out_1_iv_3\ : std_logic;
signal \uut.out_1_0_ivdup_2\ : std_logic;
signal \uut.out_1_0_iv_3\ : std_logic;
signal \uut.MAR_LD_0\ : std_logic;
signal \INVuut.out_reg.ff4.qC_net\ : std_logic;
signal \uut.g1_0\ : std_logic;
signal \uut.ir_out_m_d_3\ : std_logic;
signal \uut.AR_BUF.g0Z0Z_5\ : std_logic;
signal \uut.AR_BUF.g0_0Z0Z_0\ : std_logic;
signal \uut.ir_out_m_c_d_3\ : std_logic;
signal \uut.mar_out_2\ : std_logic;
signal \uut.mar_out_3\ : std_logic;
signal \uut.mar_out_1\ : std_logic;
signal \uut.seq.counter.T_1_fast_RNI6J9SZ0Z_3\ : std_logic;
signal \uut.D_1_3\ : std_logic;
signal \uut.seq.counter.T_1_fastZ0Z_1\ : std_logic;
signal \uut.T_3\ : std_logic;
signal \uut.un1_ROM_OE_0_cascade_\ : std_logic;
signal \uut.B_LD_0_1_tz\ : std_logic;
signal \uut.un1_ROM_OE_0\ : std_logic;
signal \uut.mem.N_7_i_m_sx_cascade_\ : std_logic;
signal \uut.B_LD_0_2_tz\ : std_logic;
signal \uut.N_7_i_m\ : std_logic;
signal \uut.AR_BUF.g0_3Z0Z_6\ : std_logic;
signal \uut.AR_BUF.g0_3Z0Z_3\ : std_logic;
signal \uut.m6\ : std_logic;
signal \uut.ROM_OE\ : std_logic;
signal \uut.mar_out_0\ : std_logic;
signal \INVuut.mar.ff4.q_neC_net\ : std_logic;
signal \uut.mar.MAR_LD_0_1\ : std_logic;
signal \_gnd_net_\ : std_logic;

signal \LED1_wire\ : std_logic;
signal \LED4_wire\ : std_logic;
signal \LED2_wire\ : std_logic;
signal \LED3_wire\ : std_logic;
signal \LED5_wire\ : std_logic;

begin
    LED1 <= \LED1_wire\;
    LED4 <= \LED4_wire\;
    LED2 <= \LED2_wire\;
    LED3 <= \LED3_wire\;
    LED5 <= \LED5_wire\;

    \LED1_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9920\,
            DIN => \N__9919\,
            DOUT => \N__9918\,
            PACKAGEPIN => \LED1_wire\
        );

    \LED1_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9920\,
            PADOUT => \N__9919\,
            PADIN => \N__9918\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3298\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED4_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9911\,
            DIN => \N__9910\,
            DOUT => \N__9909\,
            PACKAGEPIN => \LED4_wire\
        );

    \LED4_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9911\,
            PADOUT => \N__9910\,
            PADIN => \N__9909\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8161\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED2_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9902\,
            DIN => \N__9901\,
            DOUT => \N__9900\,
            PACKAGEPIN => \LED2_wire\
        );

    \LED2_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9902\,
            PADOUT => \N__9901\,
            PADIN => \N__9900\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \GNDG0\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED3_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9893\,
            DIN => \N__9892\,
            DOUT => \N__9891\,
            PACKAGEPIN => \LED3_wire\
        );

    \LED3_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9893\,
            PADOUT => \N__9892\,
            PADIN => \N__9891\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6838\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \LED5_obuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9884\,
            DIN => \N__9883\,
            DOUT => \N__9882\,
            PACKAGEPIN => \LED5_wire\
        );

    \LED5_obuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9884\,
            PADOUT => \N__9883\,
            PADIN => \N__9882\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3328\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2509\ : InMux
    port map (
            O => \N__9865\,
            I => \N__9862\
        );

    \I__2508\ : LocalMux
    port map (
            O => \N__9862\,
            I => \uut.g1_0\
        );

    \I__2507\ : InMux
    port map (
            O => \N__9859\,
            I => \N__9856\
        );

    \I__2506\ : LocalMux
    port map (
            O => \N__9856\,
            I => \N__9853\
        );

    \I__2505\ : Span4Mux_v
    port map (
            O => \N__9853\,
            I => \N__9847\
        );

    \I__2504\ : InMux
    port map (
            O => \N__9852\,
            I => \N__9844\
        );

    \I__2503\ : InMux
    port map (
            O => \N__9851\,
            I => \N__9841\
        );

    \I__2502\ : InMux
    port map (
            O => \N__9850\,
            I => \N__9837\
        );

    \I__2501\ : Span4Mux_h
    port map (
            O => \N__9847\,
            I => \N__9829\
        );

    \I__2500\ : LocalMux
    port map (
            O => \N__9844\,
            I => \N__9829\
        );

    \I__2499\ : LocalMux
    port map (
            O => \N__9841\,
            I => \N__9829\
        );

    \I__2498\ : InMux
    port map (
            O => \N__9840\,
            I => \N__9826\
        );

    \I__2497\ : LocalMux
    port map (
            O => \N__9837\,
            I => \N__9823\
        );

    \I__2496\ : InMux
    port map (
            O => \N__9836\,
            I => \N__9820\
        );

    \I__2495\ : Sp12to4
    port map (
            O => \N__9829\,
            I => \N__9815\
        );

    \I__2494\ : LocalMux
    port map (
            O => \N__9826\,
            I => \N__9815\
        );

    \I__2493\ : Odrv4
    port map (
            O => \N__9823\,
            I => \uut.ir_out_m_d_3\
        );

    \I__2492\ : LocalMux
    port map (
            O => \N__9820\,
            I => \uut.ir_out_m_d_3\
        );

    \I__2491\ : Odrv12
    port map (
            O => \N__9815\,
            I => \uut.ir_out_m_d_3\
        );

    \I__2490\ : InMux
    port map (
            O => \N__9808\,
            I => \N__9805\
        );

    \I__2489\ : LocalMux
    port map (
            O => \N__9805\,
            I => \N__9799\
        );

    \I__2488\ : InMux
    port map (
            O => \N__9804\,
            I => \N__9796\
        );

    \I__2487\ : InMux
    port map (
            O => \N__9803\,
            I => \N__9793\
        );

    \I__2486\ : InMux
    port map (
            O => \N__9802\,
            I => \N__9790\
        );

    \I__2485\ : Span4Mux_h
    port map (
            O => \N__9799\,
            I => \N__9785\
        );

    \I__2484\ : LocalMux
    port map (
            O => \N__9796\,
            I => \N__9785\
        );

    \I__2483\ : LocalMux
    port map (
            O => \N__9793\,
            I => \N__9782\
        );

    \I__2482\ : LocalMux
    port map (
            O => \N__9790\,
            I => \N__9779\
        );

    \I__2481\ : Odrv4
    port map (
            O => \N__9785\,
            I => \uut.AR_BUF.g0Z0Z_5\
        );

    \I__2480\ : Odrv12
    port map (
            O => \N__9782\,
            I => \uut.AR_BUF.g0Z0Z_5\
        );

    \I__2479\ : Odrv12
    port map (
            O => \N__9779\,
            I => \uut.AR_BUF.g0Z0Z_5\
        );

    \I__2478\ : CascadeMux
    port map (
            O => \N__9772\,
            I => \N__9768\
        );

    \I__2477\ : CascadeMux
    port map (
            O => \N__9771\,
            I => \N__9764\
        );

    \I__2476\ : InMux
    port map (
            O => \N__9768\,
            I => \N__9760\
        );

    \I__2475\ : InMux
    port map (
            O => \N__9767\,
            I => \N__9757\
        );

    \I__2474\ : InMux
    port map (
            O => \N__9764\,
            I => \N__9754\
        );

    \I__2473\ : CascadeMux
    port map (
            O => \N__9763\,
            I => \N__9751\
        );

    \I__2472\ : LocalMux
    port map (
            O => \N__9760\,
            I => \N__9748\
        );

    \I__2471\ : LocalMux
    port map (
            O => \N__9757\,
            I => \N__9743\
        );

    \I__2470\ : LocalMux
    port map (
            O => \N__9754\,
            I => \N__9743\
        );

    \I__2469\ : InMux
    port map (
            O => \N__9751\,
            I => \N__9740\
        );

    \I__2468\ : Span4Mux_s3_h
    port map (
            O => \N__9748\,
            I => \N__9736\
        );

    \I__2467\ : Span4Mux_s3_h
    port map (
            O => \N__9743\,
            I => \N__9733\
        );

    \I__2466\ : LocalMux
    port map (
            O => \N__9740\,
            I => \N__9730\
        );

    \I__2465\ : InMux
    port map (
            O => \N__9739\,
            I => \N__9727\
        );

    \I__2464\ : Odrv4
    port map (
            O => \N__9736\,
            I => \uut.AR_BUF.g0_0Z0Z_0\
        );

    \I__2463\ : Odrv4
    port map (
            O => \N__9733\,
            I => \uut.AR_BUF.g0_0Z0Z_0\
        );

    \I__2462\ : Odrv4
    port map (
            O => \N__9730\,
            I => \uut.AR_BUF.g0_0Z0Z_0\
        );

    \I__2461\ : LocalMux
    port map (
            O => \N__9727\,
            I => \uut.AR_BUF.g0_0Z0Z_0\
        );

    \I__2460\ : InMux
    port map (
            O => \N__9718\,
            I => \N__9715\
        );

    \I__2459\ : LocalMux
    port map (
            O => \N__9715\,
            I => \N__9708\
        );

    \I__2458\ : InMux
    port map (
            O => \N__9714\,
            I => \N__9705\
        );

    \I__2457\ : InMux
    port map (
            O => \N__9713\,
            I => \N__9702\
        );

    \I__2456\ : InMux
    port map (
            O => \N__9712\,
            I => \N__9697\
        );

    \I__2455\ : InMux
    port map (
            O => \N__9711\,
            I => \N__9697\
        );

    \I__2454\ : Span4Mux_v
    port map (
            O => \N__9708\,
            I => \N__9692\
        );

    \I__2453\ : LocalMux
    port map (
            O => \N__9705\,
            I => \N__9692\
        );

    \I__2452\ : LocalMux
    port map (
            O => \N__9702\,
            I => \N__9687\
        );

    \I__2451\ : LocalMux
    port map (
            O => \N__9697\,
            I => \N__9687\
        );

    \I__2450\ : Span4Mux_s3_v
    port map (
            O => \N__9692\,
            I => \N__9684\
        );

    \I__2449\ : Span12Mux_s4_h
    port map (
            O => \N__9687\,
            I => \N__9681\
        );

    \I__2448\ : Odrv4
    port map (
            O => \N__9684\,
            I => \uut.ir_out_m_c_d_3\
        );

    \I__2447\ : Odrv12
    port map (
            O => \N__9681\,
            I => \uut.ir_out_m_c_d_3\
        );

    \I__2446\ : CascadeMux
    port map (
            O => \N__9676\,
            I => \N__9672\
        );

    \I__2445\ : CascadeMux
    port map (
            O => \N__9675\,
            I => \N__9667\
        );

    \I__2444\ : InMux
    port map (
            O => \N__9672\,
            I => \N__9656\
        );

    \I__2443\ : InMux
    port map (
            O => \N__9671\,
            I => \N__9656\
        );

    \I__2442\ : InMux
    port map (
            O => \N__9670\,
            I => \N__9656\
        );

    \I__2441\ : InMux
    port map (
            O => \N__9667\,
            I => \N__9656\
        );

    \I__2440\ : InMux
    port map (
            O => \N__9666\,
            I => \N__9645\
        );

    \I__2439\ : InMux
    port map (
            O => \N__9665\,
            I => \N__9645\
        );

    \I__2438\ : LocalMux
    port map (
            O => \N__9656\,
            I => \N__9642\
        );

    \I__2437\ : InMux
    port map (
            O => \N__9655\,
            I => \N__9637\
        );

    \I__2436\ : InMux
    port map (
            O => \N__9654\,
            I => \N__9637\
        );

    \I__2435\ : InMux
    port map (
            O => \N__9653\,
            I => \N__9632\
        );

    \I__2434\ : InMux
    port map (
            O => \N__9652\,
            I => \N__9632\
        );

    \I__2433\ : InMux
    port map (
            O => \N__9651\,
            I => \N__9629\
        );

    \I__2432\ : InMux
    port map (
            O => \N__9650\,
            I => \N__9626\
        );

    \I__2431\ : LocalMux
    port map (
            O => \N__9645\,
            I => \uut.mar_out_2\
        );

    \I__2430\ : Odrv4
    port map (
            O => \N__9642\,
            I => \uut.mar_out_2\
        );

    \I__2429\ : LocalMux
    port map (
            O => \N__9637\,
            I => \uut.mar_out_2\
        );

    \I__2428\ : LocalMux
    port map (
            O => \N__9632\,
            I => \uut.mar_out_2\
        );

    \I__2427\ : LocalMux
    port map (
            O => \N__9629\,
            I => \uut.mar_out_2\
        );

    \I__2426\ : LocalMux
    port map (
            O => \N__9626\,
            I => \uut.mar_out_2\
        );

    \I__2425\ : CascadeMux
    port map (
            O => \N__9613\,
            I => \N__9604\
        );

    \I__2424\ : CascadeMux
    port map (
            O => \N__9612\,
            I => \N__9601\
        );

    \I__2423\ : CascadeMux
    port map (
            O => \N__9611\,
            I => \N__9597\
        );

    \I__2422\ : CascadeMux
    port map (
            O => \N__9610\,
            I => \N__9594\
        );

    \I__2421\ : CascadeMux
    port map (
            O => \N__9609\,
            I => \N__9591\
        );

    \I__2420\ : CascadeMux
    port map (
            O => \N__9608\,
            I => \N__9586\
        );

    \I__2419\ : InMux
    port map (
            O => \N__9607\,
            I => \N__9577\
        );

    \I__2418\ : InMux
    port map (
            O => \N__9604\,
            I => \N__9577\
        );

    \I__2417\ : InMux
    port map (
            O => \N__9601\,
            I => \N__9577\
        );

    \I__2416\ : InMux
    port map (
            O => \N__9600\,
            I => \N__9577\
        );

    \I__2415\ : InMux
    port map (
            O => \N__9597\,
            I => \N__9572\
        );

    \I__2414\ : InMux
    port map (
            O => \N__9594\,
            I => \N__9572\
        );

    \I__2413\ : InMux
    port map (
            O => \N__9591\,
            I => \N__9566\
        );

    \I__2412\ : InMux
    port map (
            O => \N__9590\,
            I => \N__9566\
        );

    \I__2411\ : InMux
    port map (
            O => \N__9589\,
            I => \N__9561\
        );

    \I__2410\ : InMux
    port map (
            O => \N__9586\,
            I => \N__9561\
        );

    \I__2409\ : LocalMux
    port map (
            O => \N__9577\,
            I => \N__9556\
        );

    \I__2408\ : LocalMux
    port map (
            O => \N__9572\,
            I => \N__9556\
        );

    \I__2407\ : InMux
    port map (
            O => \N__9571\,
            I => \N__9553\
        );

    \I__2406\ : LocalMux
    port map (
            O => \N__9566\,
            I => \uut.mar_out_3\
        );

    \I__2405\ : LocalMux
    port map (
            O => \N__9561\,
            I => \uut.mar_out_3\
        );

    \I__2404\ : Odrv4
    port map (
            O => \N__9556\,
            I => \uut.mar_out_3\
        );

    \I__2403\ : LocalMux
    port map (
            O => \N__9553\,
            I => \uut.mar_out_3\
        );

    \I__2402\ : CascadeMux
    port map (
            O => \N__9544\,
            I => \N__9540\
        );

    \I__2401\ : CascadeMux
    port map (
            O => \N__9543\,
            I => \N__9536\
        );

    \I__2400\ : InMux
    port map (
            O => \N__9540\,
            I => \N__9530\
        );

    \I__2399\ : InMux
    port map (
            O => \N__9539\,
            I => \N__9530\
        );

    \I__2398\ : InMux
    port map (
            O => \N__9536\,
            I => \N__9527\
        );

    \I__2397\ : InMux
    port map (
            O => \N__9535\,
            I => \N__9517\
        );

    \I__2396\ : LocalMux
    port map (
            O => \N__9530\,
            I => \N__9512\
        );

    \I__2395\ : LocalMux
    port map (
            O => \N__9527\,
            I => \N__9512\
        );

    \I__2394\ : InMux
    port map (
            O => \N__9526\,
            I => \N__9509\
        );

    \I__2393\ : InMux
    port map (
            O => \N__9525\,
            I => \N__9500\
        );

    \I__2392\ : InMux
    port map (
            O => \N__9524\,
            I => \N__9500\
        );

    \I__2391\ : InMux
    port map (
            O => \N__9523\,
            I => \N__9500\
        );

    \I__2390\ : InMux
    port map (
            O => \N__9522\,
            I => \N__9500\
        );

    \I__2389\ : InMux
    port map (
            O => \N__9521\,
            I => \N__9495\
        );

    \I__2388\ : InMux
    port map (
            O => \N__9520\,
            I => \N__9495\
        );

    \I__2387\ : LocalMux
    port map (
            O => \N__9517\,
            I => \N__9490\
        );

    \I__2386\ : Span4Mux_s3_v
    port map (
            O => \N__9512\,
            I => \N__9490\
        );

    \I__2385\ : LocalMux
    port map (
            O => \N__9509\,
            I => \uut.mar_out_1\
        );

    \I__2384\ : LocalMux
    port map (
            O => \N__9500\,
            I => \uut.mar_out_1\
        );

    \I__2383\ : LocalMux
    port map (
            O => \N__9495\,
            I => \uut.mar_out_1\
        );

    \I__2382\ : Odrv4
    port map (
            O => \N__9490\,
            I => \uut.mar_out_1\
        );

    \I__2381\ : InMux
    port map (
            O => \N__9481\,
            I => \N__9478\
        );

    \I__2380\ : LocalMux
    port map (
            O => \N__9478\,
            I => \N__9475\
        );

    \I__2379\ : Span4Mux_s3_h
    port map (
            O => \N__9475\,
            I => \N__9472\
        );

    \I__2378\ : Odrv4
    port map (
            O => \N__9472\,
            I => \uut.seq.counter.T_1_fast_RNI6J9SZ0Z_3\
        );

    \I__2377\ : InMux
    port map (
            O => \N__9469\,
            I => \N__9465\
        );

    \I__2376\ : InMux
    port map (
            O => \N__9468\,
            I => \N__9461\
        );

    \I__2375\ : LocalMux
    port map (
            O => \N__9465\,
            I => \N__9455\
        );

    \I__2374\ : InMux
    port map (
            O => \N__9464\,
            I => \N__9452\
        );

    \I__2373\ : LocalMux
    port map (
            O => \N__9461\,
            I => \N__9449\
        );

    \I__2372\ : InMux
    port map (
            O => \N__9460\,
            I => \N__9446\
        );

    \I__2371\ : InMux
    port map (
            O => \N__9459\,
            I => \N__9441\
        );

    \I__2370\ : InMux
    port map (
            O => \N__9458\,
            I => \N__9441\
        );

    \I__2369\ : Span4Mux_s2_v
    port map (
            O => \N__9455\,
            I => \N__9436\
        );

    \I__2368\ : LocalMux
    port map (
            O => \N__9452\,
            I => \N__9436\
        );

    \I__2367\ : Odrv12
    port map (
            O => \N__9449\,
            I => \uut.D_1_3\
        );

    \I__2366\ : LocalMux
    port map (
            O => \N__9446\,
            I => \uut.D_1_3\
        );

    \I__2365\ : LocalMux
    port map (
            O => \N__9441\,
            I => \uut.D_1_3\
        );

    \I__2364\ : Odrv4
    port map (
            O => \N__9436\,
            I => \uut.D_1_3\
        );

    \I__2363\ : InMux
    port map (
            O => \N__9427\,
            I => \N__9424\
        );

    \I__2362\ : LocalMux
    port map (
            O => \N__9424\,
            I => \N__9421\
        );

    \I__2361\ : Span4Mux_s2_h
    port map (
            O => \N__9421\,
            I => \N__9416\
        );

    \I__2360\ : InMux
    port map (
            O => \N__9420\,
            I => \N__9413\
        );

    \I__2359\ : InMux
    port map (
            O => \N__9419\,
            I => \N__9410\
        );

    \I__2358\ : Odrv4
    port map (
            O => \N__9416\,
            I => \uut.seq.counter.T_1_fastZ0Z_1\
        );

    \I__2357\ : LocalMux
    port map (
            O => \N__9413\,
            I => \uut.seq.counter.T_1_fastZ0Z_1\
        );

    \I__2356\ : LocalMux
    port map (
            O => \N__9410\,
            I => \uut.seq.counter.T_1_fastZ0Z_1\
        );

    \I__2355\ : InMux
    port map (
            O => \N__9403\,
            I => \N__9397\
        );

    \I__2354\ : InMux
    port map (
            O => \N__9402\,
            I => \N__9390\
        );

    \I__2353\ : InMux
    port map (
            O => \N__9401\,
            I => \N__9387\
        );

    \I__2352\ : InMux
    port map (
            O => \N__9400\,
            I => \N__9384\
        );

    \I__2351\ : LocalMux
    port map (
            O => \N__9397\,
            I => \N__9381\
        );

    \I__2350\ : InMux
    port map (
            O => \N__9396\,
            I => \N__9378\
        );

    \I__2349\ : InMux
    port map (
            O => \N__9395\,
            I => \N__9373\
        );

    \I__2348\ : InMux
    port map (
            O => \N__9394\,
            I => \N__9373\
        );

    \I__2347\ : InMux
    port map (
            O => \N__9393\,
            I => \N__9370\
        );

    \I__2346\ : LocalMux
    port map (
            O => \N__9390\,
            I => \N__9367\
        );

    \I__2345\ : LocalMux
    port map (
            O => \N__9387\,
            I => \N__9364\
        );

    \I__2344\ : LocalMux
    port map (
            O => \N__9384\,
            I => \N__9357\
        );

    \I__2343\ : Span4Mux_h
    port map (
            O => \N__9381\,
            I => \N__9357\
        );

    \I__2342\ : LocalMux
    port map (
            O => \N__9378\,
            I => \N__9353\
        );

    \I__2341\ : LocalMux
    port map (
            O => \N__9373\,
            I => \N__9350\
        );

    \I__2340\ : LocalMux
    port map (
            O => \N__9370\,
            I => \N__9345\
        );

    \I__2339\ : Span4Mux_h
    port map (
            O => \N__9367\,
            I => \N__9345\
        );

    \I__2338\ : Span4Mux_h
    port map (
            O => \N__9364\,
            I => \N__9342\
        );

    \I__2337\ : InMux
    port map (
            O => \N__9363\,
            I => \N__9337\
        );

    \I__2336\ : InMux
    port map (
            O => \N__9362\,
            I => \N__9337\
        );

    \I__2335\ : Span4Mux_v
    port map (
            O => \N__9357\,
            I => \N__9334\
        );

    \I__2334\ : InMux
    port map (
            O => \N__9356\,
            I => \N__9331\
        );

    \I__2333\ : Span4Mux_h
    port map (
            O => \N__9353\,
            I => \N__9324\
        );

    \I__2332\ : Span4Mux_h
    port map (
            O => \N__9350\,
            I => \N__9324\
        );

    \I__2331\ : Span4Mux_v
    port map (
            O => \N__9345\,
            I => \N__9324\
        );

    \I__2330\ : Odrv4
    port map (
            O => \N__9342\,
            I => \uut.T_3\
        );

    \I__2329\ : LocalMux
    port map (
            O => \N__9337\,
            I => \uut.T_3\
        );

    \I__2328\ : Odrv4
    port map (
            O => \N__9334\,
            I => \uut.T_3\
        );

    \I__2327\ : LocalMux
    port map (
            O => \N__9331\,
            I => \uut.T_3\
        );

    \I__2326\ : Odrv4
    port map (
            O => \N__9324\,
            I => \uut.T_3\
        );

    \I__2325\ : CascadeMux
    port map (
            O => \N__9313\,
            I => \uut.un1_ROM_OE_0_cascade_\
        );

    \I__2324\ : InMux
    port map (
            O => \N__9310\,
            I => \N__9306\
        );

    \I__2323\ : InMux
    port map (
            O => \N__9309\,
            I => \N__9303\
        );

    \I__2322\ : LocalMux
    port map (
            O => \N__9306\,
            I => \uut.B_LD_0_1_tz\
        );

    \I__2321\ : LocalMux
    port map (
            O => \N__9303\,
            I => \uut.B_LD_0_1_tz\
        );

    \I__2320\ : InMux
    port map (
            O => \N__9298\,
            I => \N__9294\
        );

    \I__2319\ : InMux
    port map (
            O => \N__9297\,
            I => \N__9291\
        );

    \I__2318\ : LocalMux
    port map (
            O => \N__9294\,
            I => \uut.un1_ROM_OE_0\
        );

    \I__2317\ : LocalMux
    port map (
            O => \N__9291\,
            I => \uut.un1_ROM_OE_0\
        );

    \I__2316\ : CascadeMux
    port map (
            O => \N__9286\,
            I => \uut.mem.N_7_i_m_sx_cascade_\
        );

    \I__2315\ : InMux
    port map (
            O => \N__9283\,
            I => \N__9280\
        );

    \I__2314\ : LocalMux
    port map (
            O => \N__9280\,
            I => \N__9275\
        );

    \I__2313\ : InMux
    port map (
            O => \N__9279\,
            I => \N__9270\
        );

    \I__2312\ : InMux
    port map (
            O => \N__9278\,
            I => \N__9270\
        );

    \I__2311\ : Span4Mux_s0_h
    port map (
            O => \N__9275\,
            I => \N__9265\
        );

    \I__2310\ : LocalMux
    port map (
            O => \N__9270\,
            I => \N__9265\
        );

    \I__2309\ : Odrv4
    port map (
            O => \N__9265\,
            I => \uut.B_LD_0_2_tz\
        );

    \I__2308\ : InMux
    port map (
            O => \N__9262\,
            I => \N__9259\
        );

    \I__2307\ : LocalMux
    port map (
            O => \N__9259\,
            I => \N__9255\
        );

    \I__2306\ : InMux
    port map (
            O => \N__9258\,
            I => \N__9252\
        );

    \I__2305\ : Span4Mux_v
    port map (
            O => \N__9255\,
            I => \N__9247\
        );

    \I__2304\ : LocalMux
    port map (
            O => \N__9252\,
            I => \N__9247\
        );

    \I__2303\ : Span4Mux_h
    port map (
            O => \N__9247\,
            I => \N__9244\
        );

    \I__2302\ : Odrv4
    port map (
            O => \N__9244\,
            I => \uut.N_7_i_m\
        );

    \I__2301\ : InMux
    port map (
            O => \N__9241\,
            I => \N__9236\
        );

    \I__2300\ : InMux
    port map (
            O => \N__9240\,
            I => \N__9233\
        );

    \I__2299\ : InMux
    port map (
            O => \N__9239\,
            I => \N__9230\
        );

    \I__2298\ : LocalMux
    port map (
            O => \N__9236\,
            I => \N__9227\
        );

    \I__2297\ : LocalMux
    port map (
            O => \N__9233\,
            I => \N__9224\
        );

    \I__2296\ : LocalMux
    port map (
            O => \N__9230\,
            I => \N__9221\
        );

    \I__2295\ : Span4Mux_s2_h
    port map (
            O => \N__9227\,
            I => \N__9217\
        );

    \I__2294\ : Span4Mux_s3_h
    port map (
            O => \N__9224\,
            I => \N__9212\
        );

    \I__2293\ : Span4Mux_h
    port map (
            O => \N__9221\,
            I => \N__9212\
        );

    \I__2292\ : InMux
    port map (
            O => \N__9220\,
            I => \N__9209\
        );

    \I__2291\ : Span4Mux_v
    port map (
            O => \N__9217\,
            I => \N__9206\
        );

    \I__2290\ : Span4Mux_v
    port map (
            O => \N__9212\,
            I => \N__9201\
        );

    \I__2289\ : LocalMux
    port map (
            O => \N__9209\,
            I => \N__9201\
        );

    \I__2288\ : Odrv4
    port map (
            O => \N__9206\,
            I => \uut.AR_BUF.g0_3Z0Z_6\
        );

    \I__2287\ : Odrv4
    port map (
            O => \N__9201\,
            I => \uut.AR_BUF.g0_3Z0Z_6\
        );

    \I__2286\ : InMux
    port map (
            O => \N__9196\,
            I => \N__9191\
        );

    \I__2285\ : CascadeMux
    port map (
            O => \N__9195\,
            I => \N__9188\
        );

    \I__2284\ : CascadeMux
    port map (
            O => \N__9194\,
            I => \N__9185\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__9191\,
            I => \N__9182\
        );

    \I__2282\ : InMux
    port map (
            O => \N__9188\,
            I => \N__9179\
        );

    \I__2281\ : InMux
    port map (
            O => \N__9185\,
            I => \N__9176\
        );

    \I__2280\ : Span4Mux_v
    port map (
            O => \N__9182\,
            I => \N__9172\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__9179\,
            I => \N__9169\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__9176\,
            I => \N__9166\
        );

    \I__2277\ : InMux
    port map (
            O => \N__9175\,
            I => \N__9163\
        );

    \I__2276\ : Span4Mux_h
    port map (
            O => \N__9172\,
            I => \N__9158\
        );

    \I__2275\ : Span4Mux_v
    port map (
            O => \N__9169\,
            I => \N__9158\
        );

    \I__2274\ : Span4Mux_v
    port map (
            O => \N__9166\,
            I => \N__9155\
        );

    \I__2273\ : LocalMux
    port map (
            O => \N__9163\,
            I => \N__9152\
        );

    \I__2272\ : Span4Mux_v
    port map (
            O => \N__9158\,
            I => \N__9147\
        );

    \I__2271\ : Span4Mux_v
    port map (
            O => \N__9155\,
            I => \N__9147\
        );

    \I__2270\ : Span4Mux_v
    port map (
            O => \N__9152\,
            I => \N__9144\
        );

    \I__2269\ : Odrv4
    port map (
            O => \N__9147\,
            I => \uut.AR_BUF.g0_3Z0Z_3\
        );

    \I__2268\ : Odrv4
    port map (
            O => \N__9144\,
            I => \uut.AR_BUF.g0_3Z0Z_3\
        );

    \I__2267\ : InMux
    port map (
            O => \N__9139\,
            I => \N__9134\
        );

    \I__2266\ : InMux
    port map (
            O => \N__9138\,
            I => \N__9130\
        );

    \I__2265\ : InMux
    port map (
            O => \N__9137\,
            I => \N__9127\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__9134\,
            I => \N__9124\
        );

    \I__2263\ : CascadeMux
    port map (
            O => \N__9133\,
            I => \N__9120\
        );

    \I__2262\ : LocalMux
    port map (
            O => \N__9130\,
            I => \N__9117\
        );

    \I__2261\ : LocalMux
    port map (
            O => \N__9127\,
            I => \N__9114\
        );

    \I__2260\ : Span4Mux_h
    port map (
            O => \N__9124\,
            I => \N__9111\
        );

    \I__2259\ : InMux
    port map (
            O => \N__9123\,
            I => \N__9107\
        );

    \I__2258\ : InMux
    port map (
            O => \N__9120\,
            I => \N__9104\
        );

    \I__2257\ : Span4Mux_h
    port map (
            O => \N__9117\,
            I => \N__9101\
        );

    \I__2256\ : Span12Mux_s2_v
    port map (
            O => \N__9114\,
            I => \N__9098\
        );

    \I__2255\ : Span4Mux_v
    port map (
            O => \N__9111\,
            I => \N__9095\
        );

    \I__2254\ : InMux
    port map (
            O => \N__9110\,
            I => \N__9092\
        );

    \I__2253\ : LocalMux
    port map (
            O => \N__9107\,
            I => \uut.m6\
        );

    \I__2252\ : LocalMux
    port map (
            O => \N__9104\,
            I => \uut.m6\
        );

    \I__2251\ : Odrv4
    port map (
            O => \N__9101\,
            I => \uut.m6\
        );

    \I__2250\ : Odrv12
    port map (
            O => \N__9098\,
            I => \uut.m6\
        );

    \I__2249\ : Odrv4
    port map (
            O => \N__9095\,
            I => \uut.m6\
        );

    \I__2248\ : LocalMux
    port map (
            O => \N__9092\,
            I => \uut.m6\
        );

    \I__2247\ : CascadeMux
    port map (
            O => \N__9079\,
            I => \N__9068\
        );

    \I__2246\ : InMux
    port map (
            O => \N__9078\,
            I => \N__9065\
        );

    \I__2245\ : InMux
    port map (
            O => \N__9077\,
            I => \N__9058\
        );

    \I__2244\ : InMux
    port map (
            O => \N__9076\,
            I => \N__9058\
        );

    \I__2243\ : InMux
    port map (
            O => \N__9075\,
            I => \N__9058\
        );

    \I__2242\ : InMux
    port map (
            O => \N__9074\,
            I => \N__9055\
        );

    \I__2241\ : InMux
    port map (
            O => \N__9073\,
            I => \N__9050\
        );

    \I__2240\ : InMux
    port map (
            O => \N__9072\,
            I => \N__9047\
        );

    \I__2239\ : CascadeMux
    port map (
            O => \N__9071\,
            I => \N__9039\
        );

    \I__2238\ : InMux
    port map (
            O => \N__9068\,
            I => \N__9034\
        );

    \I__2237\ : LocalMux
    port map (
            O => \N__9065\,
            I => \N__9029\
        );

    \I__2236\ : LocalMux
    port map (
            O => \N__9058\,
            I => \N__9026\
        );

    \I__2235\ : LocalMux
    port map (
            O => \N__9055\,
            I => \N__9023\
        );

    \I__2234\ : InMux
    port map (
            O => \N__9054\,
            I => \N__9020\
        );

    \I__2233\ : InMux
    port map (
            O => \N__9053\,
            I => \N__9017\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__9050\,
            I => \N__9012\
        );

    \I__2231\ : LocalMux
    port map (
            O => \N__9047\,
            I => \N__9012\
        );

    \I__2230\ : InMux
    port map (
            O => \N__9046\,
            I => \N__9009\
        );

    \I__2229\ : InMux
    port map (
            O => \N__9045\,
            I => \N__9006\
        );

    \I__2228\ : InMux
    port map (
            O => \N__9044\,
            I => \N__9002\
        );

    \I__2227\ : InMux
    port map (
            O => \N__9043\,
            I => \N__8995\
        );

    \I__2226\ : InMux
    port map (
            O => \N__9042\,
            I => \N__8995\
        );

    \I__2225\ : InMux
    port map (
            O => \N__9039\,
            I => \N__8995\
        );

    \I__2224\ : InMux
    port map (
            O => \N__9038\,
            I => \N__8992\
        );

    \I__2223\ : InMux
    port map (
            O => \N__9037\,
            I => \N__8989\
        );

    \I__2222\ : LocalMux
    port map (
            O => \N__9034\,
            I => \N__8986\
        );

    \I__2221\ : InMux
    port map (
            O => \N__9033\,
            I => \N__8981\
        );

    \I__2220\ : InMux
    port map (
            O => \N__9032\,
            I => \N__8978\
        );

    \I__2219\ : Span4Mux_h
    port map (
            O => \N__9029\,
            I => \N__8968\
        );

    \I__2218\ : Span4Mux_v
    port map (
            O => \N__9026\,
            I => \N__8961\
        );

    \I__2217\ : Span4Mux_v
    port map (
            O => \N__9023\,
            I => \N__8961\
        );

    \I__2216\ : LocalMux
    port map (
            O => \N__9020\,
            I => \N__8961\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__9017\,
            I => \N__8954\
        );

    \I__2214\ : Span4Mux_v
    port map (
            O => \N__9012\,
            I => \N__8954\
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__9009\,
            I => \N__8954\
        );

    \I__2212\ : LocalMux
    port map (
            O => \N__9006\,
            I => \N__8951\
        );

    \I__2211\ : InMux
    port map (
            O => \N__9005\,
            I => \N__8948\
        );

    \I__2210\ : LocalMux
    port map (
            O => \N__9002\,
            I => \N__8941\
        );

    \I__2209\ : LocalMux
    port map (
            O => \N__8995\,
            I => \N__8941\
        );

    \I__2208\ : LocalMux
    port map (
            O => \N__8992\,
            I => \N__8941\
        );

    \I__2207\ : LocalMux
    port map (
            O => \N__8989\,
            I => \N__8938\
        );

    \I__2206\ : Span4Mux_v
    port map (
            O => \N__8986\,
            I => \N__8935\
        );

    \I__2205\ : InMux
    port map (
            O => \N__8985\,
            I => \N__8932\
        );

    \I__2204\ : InMux
    port map (
            O => \N__8984\,
            I => \N__8929\
        );

    \I__2203\ : LocalMux
    port map (
            O => \N__8981\,
            I => \N__8924\
        );

    \I__2202\ : LocalMux
    port map (
            O => \N__8978\,
            I => \N__8924\
        );

    \I__2201\ : InMux
    port map (
            O => \N__8977\,
            I => \N__8920\
        );

    \I__2200\ : InMux
    port map (
            O => \N__8976\,
            I => \N__8917\
        );

    \I__2199\ : InMux
    port map (
            O => \N__8975\,
            I => \N__8908\
        );

    \I__2198\ : InMux
    port map (
            O => \N__8974\,
            I => \N__8908\
        );

    \I__2197\ : InMux
    port map (
            O => \N__8973\,
            I => \N__8908\
        );

    \I__2196\ : InMux
    port map (
            O => \N__8972\,
            I => \N__8908\
        );

    \I__2195\ : InMux
    port map (
            O => \N__8971\,
            I => \N__8905\
        );

    \I__2194\ : Sp12to4
    port map (
            O => \N__8968\,
            I => \N__8902\
        );

    \I__2193\ : Span4Mux_h
    port map (
            O => \N__8961\,
            I => \N__8897\
        );

    \I__2192\ : Span4Mux_h
    port map (
            O => \N__8954\,
            I => \N__8897\
        );

    \I__2191\ : Span12Mux_v
    port map (
            O => \N__8951\,
            I => \N__8892\
        );

    \I__2190\ : LocalMux
    port map (
            O => \N__8948\,
            I => \N__8892\
        );

    \I__2189\ : Span12Mux_s10_h
    port map (
            O => \N__8941\,
            I => \N__8889\
        );

    \I__2188\ : Span4Mux_h
    port map (
            O => \N__8938\,
            I => \N__8880\
        );

    \I__2187\ : Span4Mux_h
    port map (
            O => \N__8935\,
            I => \N__8880\
        );

    \I__2186\ : LocalMux
    port map (
            O => \N__8932\,
            I => \N__8880\
        );

    \I__2185\ : LocalMux
    port map (
            O => \N__8929\,
            I => \N__8880\
        );

    \I__2184\ : Span4Mux_s1_h
    port map (
            O => \N__8924\,
            I => \N__8877\
        );

    \I__2183\ : InMux
    port map (
            O => \N__8923\,
            I => \N__8874\
        );

    \I__2182\ : LocalMux
    port map (
            O => \N__8920\,
            I => \uut.ROM_OE\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__8917\,
            I => \uut.ROM_OE\
        );

    \I__2180\ : LocalMux
    port map (
            O => \N__8908\,
            I => \uut.ROM_OE\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__8905\,
            I => \uut.ROM_OE\
        );

    \I__2178\ : Odrv12
    port map (
            O => \N__8902\,
            I => \uut.ROM_OE\
        );

    \I__2177\ : Odrv4
    port map (
            O => \N__8897\,
            I => \uut.ROM_OE\
        );

    \I__2176\ : Odrv12
    port map (
            O => \N__8892\,
            I => \uut.ROM_OE\
        );

    \I__2175\ : Odrv12
    port map (
            O => \N__8889\,
            I => \uut.ROM_OE\
        );

    \I__2174\ : Odrv4
    port map (
            O => \N__8880\,
            I => \uut.ROM_OE\
        );

    \I__2173\ : Odrv4
    port map (
            O => \N__8877\,
            I => \uut.ROM_OE\
        );

    \I__2172\ : LocalMux
    port map (
            O => \N__8874\,
            I => \uut.ROM_OE\
        );

    \I__2171\ : InMux
    port map (
            O => \N__8851\,
            I => \N__8833\
        );

    \I__2170\ : InMux
    port map (
            O => \N__8850\,
            I => \N__8833\
        );

    \I__2169\ : InMux
    port map (
            O => \N__8849\,
            I => \N__8833\
        );

    \I__2168\ : InMux
    port map (
            O => \N__8848\,
            I => \N__8833\
        );

    \I__2167\ : InMux
    port map (
            O => \N__8847\,
            I => \N__8828\
        );

    \I__2166\ : InMux
    port map (
            O => \N__8846\,
            I => \N__8828\
        );

    \I__2165\ : InMux
    port map (
            O => \N__8845\,
            I => \N__8822\
        );

    \I__2164\ : InMux
    port map (
            O => \N__8844\,
            I => \N__8822\
        );

    \I__2163\ : InMux
    port map (
            O => \N__8843\,
            I => \N__8817\
        );

    \I__2162\ : InMux
    port map (
            O => \N__8842\,
            I => \N__8817\
        );

    \I__2161\ : LocalMux
    port map (
            O => \N__8833\,
            I => \N__8812\
        );

    \I__2160\ : LocalMux
    port map (
            O => \N__8828\,
            I => \N__8812\
        );

    \I__2159\ : InMux
    port map (
            O => \N__8827\,
            I => \N__8809\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__8822\,
            I => \uut.mar_out_0\
        );

    \I__2157\ : LocalMux
    port map (
            O => \N__8817\,
            I => \uut.mar_out_0\
        );

    \I__2156\ : Odrv4
    port map (
            O => \N__8812\,
            I => \uut.mar_out_0\
        );

    \I__2155\ : LocalMux
    port map (
            O => \N__8809\,
            I => \uut.mar_out_0\
        );

    \I__2154\ : CEMux
    port map (
            O => \N__8800\,
            I => \N__8796\
        );

    \I__2153\ : CEMux
    port map (
            O => \N__8799\,
            I => \N__8793\
        );

    \I__2152\ : LocalMux
    port map (
            O => \N__8796\,
            I => \N__8790\
        );

    \I__2151\ : LocalMux
    port map (
            O => \N__8793\,
            I => \N__8787\
        );

    \I__2150\ : Span4Mux_v
    port map (
            O => \N__8790\,
            I => \N__8784\
        );

    \I__2149\ : Span4Mux_v
    port map (
            O => \N__8787\,
            I => \N__8781\
        );

    \I__2148\ : Span4Mux_s0_v
    port map (
            O => \N__8784\,
            I => \N__8778\
        );

    \I__2147\ : Odrv4
    port map (
            O => \N__8781\,
            I => \uut.mar.MAR_LD_0_1\
        );

    \I__2146\ : Odrv4
    port map (
            O => \N__8778\,
            I => \uut.mar.MAR_LD_0_1\
        );

    \I__2145\ : CascadeMux
    port map (
            O => \N__8773\,
            I => \N__8770\
        );

    \I__2144\ : InMux
    port map (
            O => \N__8770\,
            I => \N__8762\
        );

    \I__2143\ : CascadeMux
    port map (
            O => \N__8769\,
            I => \N__8758\
        );

    \I__2142\ : InMux
    port map (
            O => \N__8768\,
            I => \N__8753\
        );

    \I__2141\ : InMux
    port map (
            O => \N__8767\,
            I => \N__8750\
        );

    \I__2140\ : InMux
    port map (
            O => \N__8766\,
            I => \N__8745\
        );

    \I__2139\ : InMux
    port map (
            O => \N__8765\,
            I => \N__8745\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__8762\,
            I => \N__8741\
        );

    \I__2137\ : InMux
    port map (
            O => \N__8761\,
            I => \N__8736\
        );

    \I__2136\ : InMux
    port map (
            O => \N__8758\,
            I => \N__8736\
        );

    \I__2135\ : InMux
    port map (
            O => \N__8757\,
            I => \N__8733\
        );

    \I__2134\ : InMux
    port map (
            O => \N__8756\,
            I => \N__8730\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__8753\,
            I => \N__8727\
        );

    \I__2132\ : LocalMux
    port map (
            O => \N__8750\,
            I => \N__8724\
        );

    \I__2131\ : LocalMux
    port map (
            O => \N__8745\,
            I => \N__8721\
        );

    \I__2130\ : InMux
    port map (
            O => \N__8744\,
            I => \N__8718\
        );

    \I__2129\ : Span4Mux_h
    port map (
            O => \N__8741\,
            I => \N__8710\
        );

    \I__2128\ : LocalMux
    port map (
            O => \N__8736\,
            I => \N__8710\
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__8733\,
            I => \N__8707\
        );

    \I__2126\ : LocalMux
    port map (
            O => \N__8730\,
            I => \N__8704\
        );

    \I__2125\ : Span4Mux_v
    port map (
            O => \N__8727\,
            I => \N__8695\
        );

    \I__2124\ : Span4Mux_v
    port map (
            O => \N__8724\,
            I => \N__8695\
        );

    \I__2123\ : Span4Mux_s0_h
    port map (
            O => \N__8721\,
            I => \N__8695\
        );

    \I__2122\ : LocalMux
    port map (
            O => \N__8718\,
            I => \N__8695\
        );

    \I__2121\ : CascadeMux
    port map (
            O => \N__8717\,
            I => \N__8692\
        );

    \I__2120\ : CascadeMux
    port map (
            O => \N__8716\,
            I => \N__8689\
        );

    \I__2119\ : InMux
    port map (
            O => \N__8715\,
            I => \N__8686\
        );

    \I__2118\ : Span4Mux_v
    port map (
            O => \N__8710\,
            I => \N__8683\
        );

    \I__2117\ : Span4Mux_v
    port map (
            O => \N__8707\,
            I => \N__8676\
        );

    \I__2116\ : Span4Mux_v
    port map (
            O => \N__8704\,
            I => \N__8676\
        );

    \I__2115\ : Span4Mux_h
    port map (
            O => \N__8695\,
            I => \N__8676\
        );

    \I__2114\ : InMux
    port map (
            O => \N__8692\,
            I => \N__8673\
        );

    \I__2113\ : InMux
    port map (
            O => \N__8689\,
            I => \N__8670\
        );

    \I__2112\ : LocalMux
    port map (
            O => \N__8686\,
            I => \uut.T_2\
        );

    \I__2111\ : Odrv4
    port map (
            O => \N__8683\,
            I => \uut.T_2\
        );

    \I__2110\ : Odrv4
    port map (
            O => \N__8676\,
            I => \uut.T_2\
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__8673\,
            I => \uut.T_2\
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__8670\,
            I => \uut.T_2\
        );

    \I__2107\ : InMux
    port map (
            O => \N__8659\,
            I => \N__8651\
        );

    \I__2106\ : InMux
    port map (
            O => \N__8658\,
            I => \N__8648\
        );

    \I__2105\ : InMux
    port map (
            O => \N__8657\,
            I => \N__8643\
        );

    \I__2104\ : InMux
    port map (
            O => \N__8656\,
            I => \N__8643\
        );

    \I__2103\ : InMux
    port map (
            O => \N__8655\,
            I => \N__8638\
        );

    \I__2102\ : InMux
    port map (
            O => \N__8654\,
            I => \N__8638\
        );

    \I__2101\ : LocalMux
    port map (
            O => \N__8651\,
            I => \N__8635\
        );

    \I__2100\ : LocalMux
    port map (
            O => \N__8648\,
            I => \N__8630\
        );

    \I__2099\ : LocalMux
    port map (
            O => \N__8643\,
            I => \N__8627\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__8638\,
            I => \N__8624\
        );

    \I__2097\ : Span12Mux_s11_h
    port map (
            O => \N__8635\,
            I => \N__8621\
        );

    \I__2096\ : InMux
    port map (
            O => \N__8634\,
            I => \N__8616\
        );

    \I__2095\ : InMux
    port map (
            O => \N__8633\,
            I => \N__8616\
        );

    \I__2094\ : Span4Mux_v
    port map (
            O => \N__8630\,
            I => \N__8611\
        );

    \I__2093\ : Span4Mux_v
    port map (
            O => \N__8627\,
            I => \N__8611\
        );

    \I__2092\ : Odrv4
    port map (
            O => \N__8624\,
            I => \uut.T_0\
        );

    \I__2091\ : Odrv12
    port map (
            O => \N__8621\,
            I => \uut.T_0\
        );

    \I__2090\ : LocalMux
    port map (
            O => \N__8616\,
            I => \uut.T_0\
        );

    \I__2089\ : Odrv4
    port map (
            O => \N__8611\,
            I => \uut.T_0\
        );

    \I__2088\ : InMux
    port map (
            O => \N__8602\,
            I => \N__8598\
        );

    \I__2087\ : CascadeMux
    port map (
            O => \N__8601\,
            I => \N__8594\
        );

    \I__2086\ : LocalMux
    port map (
            O => \N__8598\,
            I => \N__8591\
        );

    \I__2085\ : InMux
    port map (
            O => \N__8597\,
            I => \N__8586\
        );

    \I__2084\ : InMux
    port map (
            O => \N__8594\,
            I => \N__8586\
        );

    \I__2083\ : Odrv4
    port map (
            O => \N__8591\,
            I => \uut.program_counter_3\
        );

    \I__2082\ : LocalMux
    port map (
            O => \N__8586\,
            I => \uut.program_counter_3\
        );

    \I__2081\ : InMux
    port map (
            O => \N__8581\,
            I => \N__8569\
        );

    \I__2080\ : InMux
    port map (
            O => \N__8580\,
            I => \N__8569\
        );

    \I__2079\ : InMux
    port map (
            O => \N__8579\,
            I => \N__8566\
        );

    \I__2078\ : InMux
    port map (
            O => \N__8578\,
            I => \N__8559\
        );

    \I__2077\ : InMux
    port map (
            O => \N__8577\,
            I => \N__8559\
        );

    \I__2076\ : InMux
    port map (
            O => \N__8576\,
            I => \N__8559\
        );

    \I__2075\ : InMux
    port map (
            O => \N__8575\,
            I => \N__8556\
        );

    \I__2074\ : InMux
    port map (
            O => \N__8574\,
            I => \N__8553\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__8569\,
            I => \N__8546\
        );

    \I__2072\ : LocalMux
    port map (
            O => \N__8566\,
            I => \N__8541\
        );

    \I__2071\ : LocalMux
    port map (
            O => \N__8559\,
            I => \N__8541\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__8556\,
            I => \N__8536\
        );

    \I__2069\ : LocalMux
    port map (
            O => \N__8553\,
            I => \N__8536\
        );

    \I__2068\ : InMux
    port map (
            O => \N__8552\,
            I => \N__8531\
        );

    \I__2067\ : InMux
    port map (
            O => \N__8551\,
            I => \N__8531\
        );

    \I__2066\ : InMux
    port map (
            O => \N__8550\,
            I => \N__8528\
        );

    \I__2065\ : InMux
    port map (
            O => \N__8549\,
            I => \N__8525\
        );

    \I__2064\ : Span4Mux_v
    port map (
            O => \N__8546\,
            I => \N__8522\
        );

    \I__2063\ : Span4Mux_h
    port map (
            O => \N__8541\,
            I => \N__8515\
        );

    \I__2062\ : Span4Mux_s3_h
    port map (
            O => \N__8536\,
            I => \N__8515\
        );

    \I__2061\ : LocalMux
    port map (
            O => \N__8531\,
            I => \N__8515\
        );

    \I__2060\ : LocalMux
    port map (
            O => \N__8528\,
            I => \N__8510\
        );

    \I__2059\ : LocalMux
    port map (
            O => \N__8525\,
            I => \N__8510\
        );

    \I__2058\ : Odrv4
    port map (
            O => \N__8522\,
            I => \uut.D_6\
        );

    \I__2057\ : Odrv4
    port map (
            O => \N__8515\,
            I => \uut.D_6\
        );

    \I__2056\ : Odrv12
    port map (
            O => \N__8510\,
            I => \uut.D_6\
        );

    \I__2055\ : InMux
    port map (
            O => \N__8503\,
            I => \N__8500\
        );

    \I__2054\ : LocalMux
    port map (
            O => \N__8500\,
            I => \uut.program_counter_m_3\
        );

    \I__2053\ : CascadeMux
    port map (
            O => \N__8497\,
            I => \N__8492\
        );

    \I__2052\ : CascadeMux
    port map (
            O => \N__8496\,
            I => \N__8489\
        );

    \I__2051\ : InMux
    port map (
            O => \N__8495\,
            I => \N__8485\
        );

    \I__2050\ : InMux
    port map (
            O => \N__8492\,
            I => \N__8482\
        );

    \I__2049\ : InMux
    port map (
            O => \N__8489\,
            I => \N__8479\
        );

    \I__2048\ : InMux
    port map (
            O => \N__8488\,
            I => \N__8474\
        );

    \I__2047\ : LocalMux
    port map (
            O => \N__8485\,
            I => \N__8471\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__8482\,
            I => \N__8466\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__8479\,
            I => \N__8466\
        );

    \I__2044\ : CascadeMux
    port map (
            O => \N__8478\,
            I => \N__8461\
        );

    \I__2043\ : InMux
    port map (
            O => \N__8477\,
            I => \N__8458\
        );

    \I__2042\ : LocalMux
    port map (
            O => \N__8474\,
            I => \N__8455\
        );

    \I__2041\ : Span4Mux_h
    port map (
            O => \N__8471\,
            I => \N__8450\
        );

    \I__2040\ : Span4Mux_v
    port map (
            O => \N__8466\,
            I => \N__8450\
        );

    \I__2039\ : InMux
    port map (
            O => \N__8465\,
            I => \N__8445\
        );

    \I__2038\ : InMux
    port map (
            O => \N__8464\,
            I => \N__8445\
        );

    \I__2037\ : InMux
    port map (
            O => \N__8461\,
            I => \N__8442\
        );

    \I__2036\ : LocalMux
    port map (
            O => \N__8458\,
            I => \uut.acc_out_3\
        );

    \I__2035\ : Odrv12
    port map (
            O => \N__8455\,
            I => \uut.acc_out_3\
        );

    \I__2034\ : Odrv4
    port map (
            O => \N__8450\,
            I => \uut.acc_out_3\
        );

    \I__2033\ : LocalMux
    port map (
            O => \N__8445\,
            I => \uut.acc_out_3\
        );

    \I__2032\ : LocalMux
    port map (
            O => \N__8442\,
            I => \uut.acc_out_3\
        );

    \I__2031\ : CascadeMux
    port map (
            O => \N__8431\,
            I => \N__8427\
        );

    \I__2030\ : InMux
    port map (
            O => \N__8430\,
            I => \N__8423\
        );

    \I__2029\ : InMux
    port map (
            O => \N__8427\,
            I => \N__8420\
        );

    \I__2028\ : InMux
    port map (
            O => \N__8426\,
            I => \N__8417\
        );

    \I__2027\ : LocalMux
    port map (
            O => \N__8423\,
            I => \N__8411\
        );

    \I__2026\ : LocalMux
    port map (
            O => \N__8420\,
            I => \N__8411\
        );

    \I__2025\ : LocalMux
    port map (
            O => \N__8417\,
            I => \N__8408\
        );

    \I__2024\ : CascadeMux
    port map (
            O => \N__8416\,
            I => \N__8405\
        );

    \I__2023\ : Span4Mux_v
    port map (
            O => \N__8411\,
            I => \N__8401\
        );

    \I__2022\ : Span4Mux_s3_h
    port map (
            O => \N__8408\,
            I => \N__8398\
        );

    \I__2021\ : InMux
    port map (
            O => \N__8405\,
            I => \N__8393\
        );

    \I__2020\ : InMux
    port map (
            O => \N__8404\,
            I => \N__8393\
        );

    \I__2019\ : Odrv4
    port map (
            O => \N__8401\,
            I => \uut.ir_out_3\
        );

    \I__2018\ : Odrv4
    port map (
            O => \N__8398\,
            I => \uut.ir_out_3\
        );

    \I__2017\ : LocalMux
    port map (
            O => \N__8393\,
            I => \uut.ir_out_3\
        );

    \I__2016\ : InMux
    port map (
            O => \N__8386\,
            I => \N__8379\
        );

    \I__2015\ : InMux
    port map (
            O => \N__8385\,
            I => \N__8376\
        );

    \I__2014\ : InMux
    port map (
            O => \N__8384\,
            I => \N__8372\
        );

    \I__2013\ : InMux
    port map (
            O => \N__8383\,
            I => \N__8369\
        );

    \I__2012\ : InMux
    port map (
            O => \N__8382\,
            I => \N__8366\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__8379\,
            I => \N__8361\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__8376\,
            I => \N__8361\
        );

    \I__2009\ : InMux
    port map (
            O => \N__8375\,
            I => \N__8356\
        );

    \I__2008\ : LocalMux
    port map (
            O => \N__8372\,
            I => \N__8353\
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__8369\,
            I => \N__8350\
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__8366\,
            I => \N__8347\
        );

    \I__2005\ : Span4Mux_h
    port map (
            O => \N__8361\,
            I => \N__8344\
        );

    \I__2004\ : InMux
    port map (
            O => \N__8360\,
            I => \N__8341\
        );

    \I__2003\ : InMux
    port map (
            O => \N__8359\,
            I => \N__8338\
        );

    \I__2002\ : LocalMux
    port map (
            O => \N__8356\,
            I => \N__8335\
        );

    \I__2001\ : Span4Mux_s2_h
    port map (
            O => \N__8353\,
            I => \N__8332\
        );

    \I__2000\ : Span4Mux_s2_h
    port map (
            O => \N__8350\,
            I => \N__8329\
        );

    \I__1999\ : Span4Mux_s3_h
    port map (
            O => \N__8347\,
            I => \N__8324\
        );

    \I__1998\ : Span4Mux_v
    port map (
            O => \N__8344\,
            I => \N__8324\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__8341\,
            I => \N__8321\
        );

    \I__1996\ : LocalMux
    port map (
            O => \N__8338\,
            I => \uut.un5_MAR_LD\
        );

    \I__1995\ : Odrv4
    port map (
            O => \N__8335\,
            I => \uut.un5_MAR_LD\
        );

    \I__1994\ : Odrv4
    port map (
            O => \N__8332\,
            I => \uut.un5_MAR_LD\
        );

    \I__1993\ : Odrv4
    port map (
            O => \N__8329\,
            I => \uut.un5_MAR_LD\
        );

    \I__1992\ : Odrv4
    port map (
            O => \N__8324\,
            I => \uut.un5_MAR_LD\
        );

    \I__1991\ : Odrv12
    port map (
            O => \N__8321\,
            I => \uut.un5_MAR_LD\
        );

    \I__1990\ : CascadeMux
    port map (
            O => \N__8308\,
            I => \uut.AR_BUF.out_1_ivZ0Z_0_cascade_\
        );

    \I__1989\ : InMux
    port map (
            O => \N__8305\,
            I => \N__8302\
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__8302\,
            I => \N__8298\
        );

    \I__1987\ : InMux
    port map (
            O => \N__8301\,
            I => \N__8295\
        );

    \I__1986\ : Odrv4
    port map (
            O => \N__8298\,
            I => \uut.out_1_iv_2\
        );

    \I__1985\ : LocalMux
    port map (
            O => \N__8295\,
            I => \uut.out_1_iv_2\
        );

    \I__1984\ : CascadeMux
    port map (
            O => \N__8290\,
            I => \uut.out_1_iv_2_1_cascade_\
        );

    \I__1983\ : InMux
    port map (
            O => \N__8287\,
            I => \N__8283\
        );

    \I__1982\ : InMux
    port map (
            O => \N__8286\,
            I => \N__8275\
        );

    \I__1981\ : LocalMux
    port map (
            O => \N__8283\,
            I => \N__8268\
        );

    \I__1980\ : InMux
    port map (
            O => \N__8282\,
            I => \N__8265\
        );

    \I__1979\ : InMux
    port map (
            O => \N__8281\,
            I => \N__8262\
        );

    \I__1978\ : InMux
    port map (
            O => \N__8280\,
            I => \N__8257\
        );

    \I__1977\ : InMux
    port map (
            O => \N__8279\,
            I => \N__8254\
        );

    \I__1976\ : InMux
    port map (
            O => \N__8278\,
            I => \N__8250\
        );

    \I__1975\ : LocalMux
    port map (
            O => \N__8275\,
            I => \N__8247\
        );

    \I__1974\ : InMux
    port map (
            O => \N__8274\,
            I => \N__8242\
        );

    \I__1973\ : InMux
    port map (
            O => \N__8273\,
            I => \N__8242\
        );

    \I__1972\ : InMux
    port map (
            O => \N__8272\,
            I => \N__8239\
        );

    \I__1971\ : InMux
    port map (
            O => \N__8271\,
            I => \N__8236\
        );

    \I__1970\ : Span4Mux_h
    port map (
            O => \N__8268\,
            I => \N__8229\
        );

    \I__1969\ : LocalMux
    port map (
            O => \N__8265\,
            I => \N__8229\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__8262\,
            I => \N__8229\
        );

    \I__1967\ : InMux
    port map (
            O => \N__8261\,
            I => \N__8226\
        );

    \I__1966\ : InMux
    port map (
            O => \N__8260\,
            I => \N__8223\
        );

    \I__1965\ : LocalMux
    port map (
            O => \N__8257\,
            I => \N__8218\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__8254\,
            I => \N__8218\
        );

    \I__1963\ : InMux
    port map (
            O => \N__8253\,
            I => \N__8215\
        );

    \I__1962\ : LocalMux
    port map (
            O => \N__8250\,
            I => \N__8210\
        );

    \I__1961\ : Span4Mux_v
    port map (
            O => \N__8247\,
            I => \N__8210\
        );

    \I__1960\ : LocalMux
    port map (
            O => \N__8242\,
            I => \N__8205\
        );

    \I__1959\ : LocalMux
    port map (
            O => \N__8239\,
            I => \N__8205\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__8236\,
            I => \N__8200\
        );

    \I__1957\ : Span4Mux_v
    port map (
            O => \N__8229\,
            I => \N__8200\
        );

    \I__1956\ : LocalMux
    port map (
            O => \N__8226\,
            I => \N__8197\
        );

    \I__1955\ : LocalMux
    port map (
            O => \N__8223\,
            I => \N__8194\
        );

    \I__1954\ : Span4Mux_v
    port map (
            O => \N__8218\,
            I => \N__8191\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__8215\,
            I => \N__8188\
        );

    \I__1952\ : Span4Mux_v
    port map (
            O => \N__8210\,
            I => \N__8183\
        );

    \I__1951\ : Span4Mux_h
    port map (
            O => \N__8205\,
            I => \N__8183\
        );

    \I__1950\ : Span4Mux_h
    port map (
            O => \N__8200\,
            I => \N__8178\
        );

    \I__1949\ : Span4Mux_s2_h
    port map (
            O => \N__8197\,
            I => \N__8178\
        );

    \I__1948\ : Span12Mux_s8_h
    port map (
            O => \N__8194\,
            I => \N__8175\
        );

    \I__1947\ : Sp12to4
    port map (
            O => \N__8191\,
            I => \N__8170\
        );

    \I__1946\ : Span12Mux_v
    port map (
            O => \N__8188\,
            I => \N__8170\
        );

    \I__1945\ : Odrv4
    port map (
            O => \N__8183\,
            I => \uut.OUT_LD\
        );

    \I__1944\ : Odrv4
    port map (
            O => \N__8178\,
            I => \uut.OUT_LD\
        );

    \I__1943\ : Odrv12
    port map (
            O => \N__8175\,
            I => \uut.OUT_LD\
        );

    \I__1942\ : Odrv12
    port map (
            O => \N__8170\,
            I => \uut.OUT_LD\
        );

    \I__1941\ : IoInMux
    port map (
            O => \N__8161\,
            I => \N__8158\
        );

    \I__1940\ : LocalMux
    port map (
            O => \N__8158\,
            I => \N__8154\
        );

    \I__1939\ : InMux
    port map (
            O => \N__8157\,
            I => \N__8151\
        );

    \I__1938\ : Span12Mux_s0_h
    port map (
            O => \N__8154\,
            I => \N__8148\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__8151\,
            I => \N__8145\
        );

    \I__1936\ : Odrv12
    port map (
            O => \N__8148\,
            I => \LED4_c\
        );

    \I__1935\ : Odrv4
    port map (
            O => \N__8145\,
            I => \LED4_c\
        );

    \I__1934\ : InMux
    port map (
            O => \N__8140\,
            I => \N__8137\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__8137\,
            I => \uut.alu_out_m_3\
        );

    \I__1932\ : CascadeMux
    port map (
            O => \N__8134\,
            I => \uut.m15_cascade_\
        );

    \I__1931\ : InMux
    port map (
            O => \N__8131\,
            I => \N__8128\
        );

    \I__1930\ : LocalMux
    port map (
            O => \N__8128\,
            I => \uut.out_1_iv_3\
        );

    \I__1929\ : CascadeMux
    port map (
            O => \N__8125\,
            I => \N__8122\
        );

    \I__1928\ : InMux
    port map (
            O => \N__8122\,
            I => \N__8118\
        );

    \I__1927\ : InMux
    port map (
            O => \N__8121\,
            I => \N__8115\
        );

    \I__1926\ : LocalMux
    port map (
            O => \N__8118\,
            I => \N__8112\
        );

    \I__1925\ : LocalMux
    port map (
            O => \N__8115\,
            I => \N__8109\
        );

    \I__1924\ : Span4Mux_s3_v
    port map (
            O => \N__8112\,
            I => \N__8103\
        );

    \I__1923\ : Span4Mux_s0_h
    port map (
            O => \N__8109\,
            I => \N__8103\
        );

    \I__1922\ : InMux
    port map (
            O => \N__8108\,
            I => \N__8100\
        );

    \I__1921\ : Span4Mux_h
    port map (
            O => \N__8103\,
            I => \N__8095\
        );

    \I__1920\ : LocalMux
    port map (
            O => \N__8100\,
            I => \N__8092\
        );

    \I__1919\ : InMux
    port map (
            O => \N__8099\,
            I => \N__8089\
        );

    \I__1918\ : InMux
    port map (
            O => \N__8098\,
            I => \N__8086\
        );

    \I__1917\ : Odrv4
    port map (
            O => \N__8095\,
            I => \uut.out_1_0_ivdup_2\
        );

    \I__1916\ : Odrv12
    port map (
            O => \N__8092\,
            I => \uut.out_1_0_ivdup_2\
        );

    \I__1915\ : LocalMux
    port map (
            O => \N__8089\,
            I => \uut.out_1_0_ivdup_2\
        );

    \I__1914\ : LocalMux
    port map (
            O => \N__8086\,
            I => \uut.out_1_0_ivdup_2\
        );

    \I__1913\ : InMux
    port map (
            O => \N__8077\,
            I => \N__8074\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__8074\,
            I => \N__8070\
        );

    \I__1911\ : InMux
    port map (
            O => \N__8073\,
            I => \N__8067\
        );

    \I__1910\ : Span4Mux_s3_v
    port map (
            O => \N__8070\,
            I => \N__8063\
        );

    \I__1909\ : LocalMux
    port map (
            O => \N__8067\,
            I => \N__8060\
        );

    \I__1908\ : InMux
    port map (
            O => \N__8066\,
            I => \N__8057\
        );

    \I__1907\ : Span4Mux_h
    port map (
            O => \N__8063\,
            I => \N__8050\
        );

    \I__1906\ : Span4Mux_s3_v
    port map (
            O => \N__8060\,
            I => \N__8050\
        );

    \I__1905\ : LocalMux
    port map (
            O => \N__8057\,
            I => \N__8050\
        );

    \I__1904\ : Odrv4
    port map (
            O => \N__8050\,
            I => \uut.out_1_0_iv_3\
        );

    \I__1903\ : CascadeMux
    port map (
            O => \N__8047\,
            I => \N__8044\
        );

    \I__1902\ : InMux
    port map (
            O => \N__8044\,
            I => \N__8038\
        );

    \I__1901\ : InMux
    port map (
            O => \N__8043\,
            I => \N__8038\
        );

    \I__1900\ : LocalMux
    port map (
            O => \N__8038\,
            I => \N__8035\
        );

    \I__1899\ : Odrv12
    port map (
            O => \N__8035\,
            I => \uut.MAR_LD_0\
        );

    \I__1898\ : InMux
    port map (
            O => \N__8032\,
            I => \N__8028\
        );

    \I__1897\ : CEMux
    port map (
            O => \N__8031\,
            I => \N__8024\
        );

    \I__1896\ : LocalMux
    port map (
            O => \N__8028\,
            I => \N__8020\
        );

    \I__1895\ : CEMux
    port map (
            O => \N__8027\,
            I => \N__8017\
        );

    \I__1894\ : LocalMux
    port map (
            O => \N__8024\,
            I => \N__8014\
        );

    \I__1893\ : InMux
    port map (
            O => \N__8023\,
            I => \N__8011\
        );

    \I__1892\ : Span4Mux_h
    port map (
            O => \N__8020\,
            I => \N__8008\
        );

    \I__1891\ : LocalMux
    port map (
            O => \N__8017\,
            I => \N__8005\
        );

    \I__1890\ : Span4Mux_s0_h
    port map (
            O => \N__8014\,
            I => \N__8002\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__8011\,
            I => \N__7999\
        );

    \I__1888\ : Span4Mux_h
    port map (
            O => \N__8008\,
            I => \N__7996\
        );

    \I__1887\ : Odrv12
    port map (
            O => \N__8005\,
            I => \uut.AR_LD\
        );

    \I__1886\ : Odrv4
    port map (
            O => \N__8002\,
            I => \uut.AR_LD\
        );

    \I__1885\ : Odrv4
    port map (
            O => \N__7999\,
            I => \uut.AR_LD\
        );

    \I__1884\ : Odrv4
    port map (
            O => \N__7996\,
            I => \uut.AR_LD\
        );

    \I__1883\ : InMux
    port map (
            O => \N__7987\,
            I => \N__7982\
        );

    \I__1882\ : InMux
    port map (
            O => \N__7986\,
            I => \N__7979\
        );

    \I__1881\ : InMux
    port map (
            O => \N__7985\,
            I => \N__7976\
        );

    \I__1880\ : LocalMux
    port map (
            O => \N__7982\,
            I => \N__7971\
        );

    \I__1879\ : LocalMux
    port map (
            O => \N__7979\,
            I => \N__7966\
        );

    \I__1878\ : LocalMux
    port map (
            O => \N__7976\,
            I => \N__7966\
        );

    \I__1877\ : CascadeMux
    port map (
            O => \N__7975\,
            I => \N__7962\
        );

    \I__1876\ : InMux
    port map (
            O => \N__7974\,
            I => \N__7959\
        );

    \I__1875\ : Span4Mux_v
    port map (
            O => \N__7971\,
            I => \N__7954\
        );

    \I__1874\ : Span4Mux_v
    port map (
            O => \N__7966\,
            I => \N__7954\
        );

    \I__1873\ : InMux
    port map (
            O => \N__7965\,
            I => \N__7949\
        );

    \I__1872\ : InMux
    port map (
            O => \N__7962\,
            I => \N__7949\
        );

    \I__1871\ : LocalMux
    port map (
            O => \N__7959\,
            I => \N__7946\
        );

    \I__1870\ : Odrv4
    port map (
            O => \N__7954\,
            I => \uut.un14_MAR_LD\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__7949\,
            I => \uut.un14_MAR_LD\
        );

    \I__1868\ : Odrv4
    port map (
            O => \N__7946\,
            I => \uut.un14_MAR_LD\
        );

    \I__1867\ : InMux
    port map (
            O => \N__7939\,
            I => \N__7936\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__7936\,
            I => \N__7930\
        );

    \I__1865\ : InMux
    port map (
            O => \N__7935\,
            I => \N__7926\
        );

    \I__1864\ : InMux
    port map (
            O => \N__7934\,
            I => \N__7921\
        );

    \I__1863\ : InMux
    port map (
            O => \N__7933\,
            I => \N__7921\
        );

    \I__1862\ : Span4Mux_s1_h
    port map (
            O => \N__7930\,
            I => \N__7918\
        );

    \I__1861\ : InMux
    port map (
            O => \N__7929\,
            I => \N__7915\
        );

    \I__1860\ : LocalMux
    port map (
            O => \N__7926\,
            I => \N__7912\
        );

    \I__1859\ : LocalMux
    port map (
            O => \N__7921\,
            I => \N__7909\
        );

    \I__1858\ : Span4Mux_v
    port map (
            O => \N__7918\,
            I => \N__7904\
        );

    \I__1857\ : LocalMux
    port map (
            O => \N__7915\,
            I => \N__7904\
        );

    \I__1856\ : Span4Mux_s3_h
    port map (
            O => \N__7912\,
            I => \N__7899\
        );

    \I__1855\ : Span4Mux_h
    port map (
            O => \N__7909\,
            I => \N__7899\
        );

    \I__1854\ : Odrv4
    port map (
            O => \N__7904\,
            I => \uut.un8_MAR_LD\
        );

    \I__1853\ : Odrv4
    port map (
            O => \N__7899\,
            I => \uut.un8_MAR_LD\
        );

    \I__1852\ : InMux
    port map (
            O => \N__7894\,
            I => \N__7889\
        );

    \I__1851\ : InMux
    port map (
            O => \N__7893\,
            I => \N__7886\
        );

    \I__1850\ : InMux
    port map (
            O => \N__7892\,
            I => \N__7883\
        );

    \I__1849\ : LocalMux
    port map (
            O => \N__7889\,
            I => \N__7880\
        );

    \I__1848\ : LocalMux
    port map (
            O => \N__7886\,
            I => \N__7877\
        );

    \I__1847\ : LocalMux
    port map (
            O => \N__7883\,
            I => \N__7874\
        );

    \I__1846\ : Span4Mux_s3_v
    port map (
            O => \N__7880\,
            I => \N__7869\
        );

    \I__1845\ : Span4Mux_v
    port map (
            O => \N__7877\,
            I => \N__7864\
        );

    \I__1844\ : Span4Mux_s3_h
    port map (
            O => \N__7874\,
            I => \N__7864\
        );

    \I__1843\ : InMux
    port map (
            O => \N__7873\,
            I => \N__7859\
        );

    \I__1842\ : InMux
    port map (
            O => \N__7872\,
            I => \N__7859\
        );

    \I__1841\ : Odrv4
    port map (
            O => \N__7869\,
            I => \uut.un1_IR_OE_4_1\
        );

    \I__1840\ : Odrv4
    port map (
            O => \N__7864\,
            I => \uut.un1_IR_OE_4_1\
        );

    \I__1839\ : LocalMux
    port map (
            O => \N__7859\,
            I => \uut.un1_IR_OE_4_1\
        );

    \I__1838\ : InMux
    port map (
            O => \N__7852\,
            I => \N__7849\
        );

    \I__1837\ : LocalMux
    port map (
            O => \N__7849\,
            I => \uut.pc.un1_inc_0_0\
        );

    \I__1836\ : CascadeMux
    port map (
            O => \N__7846\,
            I => \uut.ir_out_m_d_3_cascade_\
        );

    \I__1835\ : InMux
    port map (
            O => \N__7843\,
            I => \N__7840\
        );

    \I__1834\ : LocalMux
    port map (
            O => \N__7840\,
            I => \uut.pc.g0_sn\
        );

    \I__1833\ : InMux
    port map (
            O => \N__7837\,
            I => \N__7833\
        );

    \I__1832\ : InMux
    port map (
            O => \N__7836\,
            I => \N__7830\
        );

    \I__1831\ : LocalMux
    port map (
            O => \N__7833\,
            I => \N__7827\
        );

    \I__1830\ : LocalMux
    port map (
            O => \N__7830\,
            I => \N__7824\
        );

    \I__1829\ : Span12Mux_s10_h
    port map (
            O => \N__7827\,
            I => \N__7821\
        );

    \I__1828\ : Span4Mux_v
    port map (
            O => \N__7824\,
            I => \N__7818\
        );

    \I__1827\ : Odrv12
    port map (
            O => \N__7821\,
            I => \uut.seq.counter.T_1Z0Z_4\
        );

    \I__1826\ : Odrv4
    port map (
            O => \N__7818\,
            I => \uut.seq.counter.T_1Z0Z_4\
        );

    \I__1825\ : CascadeMux
    port map (
            O => \N__7813\,
            I => \uut.AR_BUF.out_1_ivdupZ0Z_0_cascade_\
        );

    \I__1824\ : InMux
    port map (
            O => \N__7810\,
            I => \N__7807\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__7807\,
            I => \uut.g0_0\
        );

    \I__1822\ : InMux
    port map (
            O => \N__7804\,
            I => \N__7800\
        );

    \I__1821\ : CascadeMux
    port map (
            O => \N__7803\,
            I => \N__7797\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__7800\,
            I => \N__7794\
        );

    \I__1819\ : InMux
    port map (
            O => \N__7797\,
            I => \N__7791\
        );

    \I__1818\ : Odrv4
    port map (
            O => \N__7794\,
            I => \uut.AR_out_3\
        );

    \I__1817\ : LocalMux
    port map (
            O => \N__7791\,
            I => \uut.AR_out_3\
        );

    \I__1816\ : CascadeMux
    port map (
            O => \N__7786\,
            I => \uut.g1_cascade_\
        );

    \I__1815\ : InMux
    port map (
            O => \N__7783\,
            I => \N__7776\
        );

    \I__1814\ : InMux
    port map (
            O => \N__7782\,
            I => \N__7773\
        );

    \I__1813\ : InMux
    port map (
            O => \N__7781\,
            I => \N__7770\
        );

    \I__1812\ : InMux
    port map (
            O => \N__7780\,
            I => \N__7765\
        );

    \I__1811\ : InMux
    port map (
            O => \N__7779\,
            I => \N__7765\
        );

    \I__1810\ : LocalMux
    port map (
            O => \N__7776\,
            I => \N__7755\
        );

    \I__1809\ : LocalMux
    port map (
            O => \N__7773\,
            I => \N__7748\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__7770\,
            I => \N__7748\
        );

    \I__1807\ : LocalMux
    port map (
            O => \N__7765\,
            I => \N__7748\
        );

    \I__1806\ : InMux
    port map (
            O => \N__7764\,
            I => \N__7745\
        );

    \I__1805\ : InMux
    port map (
            O => \N__7763\,
            I => \N__7742\
        );

    \I__1804\ : InMux
    port map (
            O => \N__7762\,
            I => \N__7739\
        );

    \I__1803\ : InMux
    port map (
            O => \N__7761\,
            I => \N__7736\
        );

    \I__1802\ : InMux
    port map (
            O => \N__7760\,
            I => \N__7733\
        );

    \I__1801\ : InMux
    port map (
            O => \N__7759\,
            I => \N__7728\
        );

    \I__1800\ : InMux
    port map (
            O => \N__7758\,
            I => \N__7728\
        );

    \I__1799\ : Span4Mux_v
    port map (
            O => \N__7755\,
            I => \N__7725\
        );

    \I__1798\ : Span4Mux_v
    port map (
            O => \N__7748\,
            I => \N__7722\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__7745\,
            I => \N__7715\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__7742\,
            I => \N__7715\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__7739\,
            I => \N__7715\
        );

    \I__1794\ : LocalMux
    port map (
            O => \N__7736\,
            I => \N__7708\
        );

    \I__1793\ : LocalMux
    port map (
            O => \N__7733\,
            I => \N__7708\
        );

    \I__1792\ : LocalMux
    port map (
            O => \N__7728\,
            I => \N__7708\
        );

    \I__1791\ : Odrv4
    port map (
            O => \N__7725\,
            I => \uut.T_2_rep1_RNI6BLF1\
        );

    \I__1790\ : Odrv4
    port map (
            O => \N__7722\,
            I => \uut.T_2_rep1_RNI6BLF1\
        );

    \I__1789\ : Odrv4
    port map (
            O => \N__7715\,
            I => \uut.T_2_rep1_RNI6BLF1\
        );

    \I__1788\ : Odrv4
    port map (
            O => \N__7708\,
            I => \uut.T_2_rep1_RNI6BLF1\
        );

    \I__1787\ : InMux
    port map (
            O => \N__7699\,
            I => \N__7696\
        );

    \I__1786\ : LocalMux
    port map (
            O => \N__7696\,
            I => \uut.AR_BUF.g0_1_0\
        );

    \I__1785\ : InMux
    port map (
            O => \N__7693\,
            I => \N__7689\
        );

    \I__1784\ : InMux
    port map (
            O => \N__7692\,
            I => \N__7685\
        );

    \I__1783\ : LocalMux
    port map (
            O => \N__7689\,
            I => \N__7681\
        );

    \I__1782\ : InMux
    port map (
            O => \N__7688\,
            I => \N__7677\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__7685\,
            I => \N__7674\
        );

    \I__1780\ : InMux
    port map (
            O => \N__7684\,
            I => \N__7671\
        );

    \I__1779\ : Span4Mux_h
    port map (
            O => \N__7681\,
            I => \N__7668\
        );

    \I__1778\ : InMux
    port map (
            O => \N__7680\,
            I => \N__7665\
        );

    \I__1777\ : LocalMux
    port map (
            O => \N__7677\,
            I => \N__7662\
        );

    \I__1776\ : Span12Mux_s7_v
    port map (
            O => \N__7674\,
            I => \N__7657\
        );

    \I__1775\ : LocalMux
    port map (
            O => \N__7671\,
            I => \N__7657\
        );

    \I__1774\ : Span4Mux_v
    port map (
            O => \N__7668\,
            I => \N__7652\
        );

    \I__1773\ : LocalMux
    port map (
            O => \N__7665\,
            I => \N__7652\
        );

    \I__1772\ : Odrv12
    port map (
            O => \N__7662\,
            I => \uut.alu_out_m_1\
        );

    \I__1771\ : Odrv12
    port map (
            O => \N__7657\,
            I => \uut.alu_out_m_1\
        );

    \I__1770\ : Odrv4
    port map (
            O => \N__7652\,
            I => \uut.alu_out_m_1\
        );

    \I__1769\ : InMux
    port map (
            O => \N__7645\,
            I => \N__7640\
        );

    \I__1768\ : InMux
    port map (
            O => \N__7644\,
            I => \N__7637\
        );

    \I__1767\ : InMux
    port map (
            O => \N__7643\,
            I => \N__7633\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__7640\,
            I => \N__7630\
        );

    \I__1765\ : LocalMux
    port map (
            O => \N__7637\,
            I => \N__7627\
        );

    \I__1764\ : InMux
    port map (
            O => \N__7636\,
            I => \N__7624\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__7633\,
            I => \N__7620\
        );

    \I__1762\ : Span4Mux_s2_v
    port map (
            O => \N__7630\,
            I => \N__7617\
        );

    \I__1761\ : Span12Mux_s10_h
    port map (
            O => \N__7627\,
            I => \N__7612\
        );

    \I__1760\ : LocalMux
    port map (
            O => \N__7624\,
            I => \N__7612\
        );

    \I__1759\ : InMux
    port map (
            O => \N__7623\,
            I => \N__7609\
        );

    \I__1758\ : Span12Mux_v
    port map (
            O => \N__7620\,
            I => \N__7606\
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__7617\,
            I => \uut.N_11_i_m\
        );

    \I__1756\ : Odrv12
    port map (
            O => \N__7612\,
            I => \uut.N_11_i_m\
        );

    \I__1755\ : LocalMux
    port map (
            O => \N__7609\,
            I => \uut.N_11_i_m\
        );

    \I__1754\ : Odrv12
    port map (
            O => \N__7606\,
            I => \uut.N_11_i_m\
        );

    \I__1753\ : InMux
    port map (
            O => \N__7597\,
            I => \N__7593\
        );

    \I__1752\ : InMux
    port map (
            O => \N__7596\,
            I => \N__7590\
        );

    \I__1751\ : LocalMux
    port map (
            O => \N__7593\,
            I => \N__7586\
        );

    \I__1750\ : LocalMux
    port map (
            O => \N__7590\,
            I => \N__7583\
        );

    \I__1749\ : InMux
    port map (
            O => \N__7589\,
            I => \N__7580\
        );

    \I__1748\ : Span4Mux_s3_v
    port map (
            O => \N__7586\,
            I => \N__7576\
        );

    \I__1747\ : Span4Mux_s3_v
    port map (
            O => \N__7583\,
            I => \N__7571\
        );

    \I__1746\ : LocalMux
    port map (
            O => \N__7580\,
            I => \N__7571\
        );

    \I__1745\ : InMux
    port map (
            O => \N__7579\,
            I => \N__7568\
        );

    \I__1744\ : Span4Mux_v
    port map (
            O => \N__7576\,
            I => \N__7562\
        );

    \I__1743\ : Span4Mux_v
    port map (
            O => \N__7571\,
            I => \N__7562\
        );

    \I__1742\ : LocalMux
    port map (
            O => \N__7568\,
            I => \N__7559\
        );

    \I__1741\ : InMux
    port map (
            O => \N__7567\,
            I => \N__7556\
        );

    \I__1740\ : Odrv4
    port map (
            O => \N__7562\,
            I => \uut.out_1_1_iv_3dup_1\
        );

    \I__1739\ : Odrv4
    port map (
            O => \N__7559\,
            I => \uut.out_1_1_iv_3dup_1\
        );

    \I__1738\ : LocalMux
    port map (
            O => \N__7556\,
            I => \uut.out_1_1_iv_3dup_1\
        );

    \I__1737\ : InMux
    port map (
            O => \N__7549\,
            I => \N__7544\
        );

    \I__1736\ : InMux
    port map (
            O => \N__7548\,
            I => \N__7541\
        );

    \I__1735\ : InMux
    port map (
            O => \N__7547\,
            I => \N__7538\
        );

    \I__1734\ : LocalMux
    port map (
            O => \N__7544\,
            I => \N__7535\
        );

    \I__1733\ : LocalMux
    port map (
            O => \N__7541\,
            I => \N__7532\
        );

    \I__1732\ : LocalMux
    port map (
            O => \N__7538\,
            I => \N__7529\
        );

    \I__1731\ : Span4Mux_h
    port map (
            O => \N__7535\,
            I => \N__7526\
        );

    \I__1730\ : Span4Mux_h
    port map (
            O => \N__7532\,
            I => \N__7523\
        );

    \I__1729\ : Odrv12
    port map (
            O => \N__7529\,
            I => \uut.b_reg_out_1\
        );

    \I__1728\ : Odrv4
    port map (
            O => \N__7526\,
            I => \uut.b_reg_out_1\
        );

    \I__1727\ : Odrv4
    port map (
            O => \N__7523\,
            I => \uut.b_reg_out_1\
        );

    \I__1726\ : CEMux
    port map (
            O => \N__7516\,
            I => \N__7511\
        );

    \I__1725\ : CEMux
    port map (
            O => \N__7515\,
            I => \N__7507\
        );

    \I__1724\ : CEMux
    port map (
            O => \N__7514\,
            I => \N__7504\
        );

    \I__1723\ : LocalMux
    port map (
            O => \N__7511\,
            I => \N__7500\
        );

    \I__1722\ : CEMux
    port map (
            O => \N__7510\,
            I => \N__7497\
        );

    \I__1721\ : LocalMux
    port map (
            O => \N__7507\,
            I => \N__7494\
        );

    \I__1720\ : LocalMux
    port map (
            O => \N__7504\,
            I => \N__7491\
        );

    \I__1719\ : CEMux
    port map (
            O => \N__7503\,
            I => \N__7488\
        );

    \I__1718\ : Span4Mux_h
    port map (
            O => \N__7500\,
            I => \N__7482\
        );

    \I__1717\ : LocalMux
    port map (
            O => \N__7497\,
            I => \N__7482\
        );

    \I__1716\ : Span4Mux_v
    port map (
            O => \N__7494\,
            I => \N__7476\
        );

    \I__1715\ : Span4Mux_v
    port map (
            O => \N__7491\,
            I => \N__7476\
        );

    \I__1714\ : LocalMux
    port map (
            O => \N__7488\,
            I => \N__7473\
        );

    \I__1713\ : CEMux
    port map (
            O => \N__7487\,
            I => \N__7470\
        );

    \I__1712\ : Span4Mux_v
    port map (
            O => \N__7482\,
            I => \N__7467\
        );

    \I__1711\ : CEMux
    port map (
            O => \N__7481\,
            I => \N__7464\
        );

    \I__1710\ : Span4Mux_s2_v
    port map (
            O => \N__7476\,
            I => \N__7461\
        );

    \I__1709\ : Span4Mux_v
    port map (
            O => \N__7473\,
            I => \N__7458\
        );

    \I__1708\ : LocalMux
    port map (
            O => \N__7470\,
            I => \N__7455\
        );

    \I__1707\ : Span4Mux_h
    port map (
            O => \N__7467\,
            I => \N__7450\
        );

    \I__1706\ : LocalMux
    port map (
            O => \N__7464\,
            I => \N__7450\
        );

    \I__1705\ : Span4Mux_h
    port map (
            O => \N__7461\,
            I => \N__7447\
        );

    \I__1704\ : Span4Mux_h
    port map (
            O => \N__7458\,
            I => \N__7444\
        );

    \I__1703\ : Span4Mux_h
    port map (
            O => \N__7455\,
            I => \N__7439\
        );

    \I__1702\ : Span4Mux_s1_h
    port map (
            O => \N__7450\,
            I => \N__7439\
        );

    \I__1701\ : Odrv4
    port map (
            O => \N__7447\,
            I => \uut.B_LD_0_i\
        );

    \I__1700\ : Odrv4
    port map (
            O => \N__7444\,
            I => \uut.B_LD_0_i\
        );

    \I__1699\ : Odrv4
    port map (
            O => \N__7439\,
            I => \uut.B_LD_0_i\
        );

    \I__1698\ : CEMux
    port map (
            O => \N__7432\,
            I => \N__7429\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__7429\,
            I => \N__7425\
        );

    \I__1696\ : CEMux
    port map (
            O => \N__7428\,
            I => \N__7422\
        );

    \I__1695\ : Span4Mux_s2_v
    port map (
            O => \N__7425\,
            I => \N__7407\
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__7422\,
            I => \N__7407\
        );

    \I__1693\ : InMux
    port map (
            O => \N__7421\,
            I => \N__7392\
        );

    \I__1692\ : InMux
    port map (
            O => \N__7420\,
            I => \N__7392\
        );

    \I__1691\ : InMux
    port map (
            O => \N__7419\,
            I => \N__7392\
        );

    \I__1690\ : InMux
    port map (
            O => \N__7418\,
            I => \N__7392\
        );

    \I__1689\ : InMux
    port map (
            O => \N__7417\,
            I => \N__7387\
        );

    \I__1688\ : InMux
    port map (
            O => \N__7416\,
            I => \N__7387\
        );

    \I__1687\ : InMux
    port map (
            O => \N__7415\,
            I => \N__7383\
        );

    \I__1686\ : InMux
    port map (
            O => \N__7414\,
            I => \N__7378\
        );

    \I__1685\ : InMux
    port map (
            O => \N__7413\,
            I => \N__7378\
        );

    \I__1684\ : InMux
    port map (
            O => \N__7412\,
            I => \N__7375\
        );

    \I__1683\ : Span4Mux_v
    port map (
            O => \N__7407\,
            I => \N__7372\
        );

    \I__1682\ : InMux
    port map (
            O => \N__7406\,
            I => \N__7369\
        );

    \I__1681\ : InMux
    port map (
            O => \N__7405\,
            I => \N__7364\
        );

    \I__1680\ : InMux
    port map (
            O => \N__7404\,
            I => \N__7364\
        );

    \I__1679\ : InMux
    port map (
            O => \N__7403\,
            I => \N__7361\
        );

    \I__1678\ : InMux
    port map (
            O => \N__7402\,
            I => \N__7357\
        );

    \I__1677\ : CEMux
    port map (
            O => \N__7401\,
            I => \N__7354\
        );

    \I__1676\ : LocalMux
    port map (
            O => \N__7392\,
            I => \N__7351\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__7387\,
            I => \N__7348\
        );

    \I__1674\ : InMux
    port map (
            O => \N__7386\,
            I => \N__7345\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__7383\,
            I => \N__7340\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__7378\,
            I => \N__7340\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__7375\,
            I => \N__7329\
        );

    \I__1670\ : Span4Mux_h
    port map (
            O => \N__7372\,
            I => \N__7329\
        );

    \I__1669\ : LocalMux
    port map (
            O => \N__7369\,
            I => \N__7329\
        );

    \I__1668\ : LocalMux
    port map (
            O => \N__7364\,
            I => \N__7329\
        );

    \I__1667\ : LocalMux
    port map (
            O => \N__7361\,
            I => \N__7329\
        );

    \I__1666\ : CascadeMux
    port map (
            O => \N__7360\,
            I => \N__7324\
        );

    \I__1665\ : LocalMux
    port map (
            O => \N__7357\,
            I => \N__7321\
        );

    \I__1664\ : LocalMux
    port map (
            O => \N__7354\,
            I => \N__7312\
        );

    \I__1663\ : Span4Mux_s2_v
    port map (
            O => \N__7351\,
            I => \N__7312\
        );

    \I__1662\ : Span4Mux_s2_v
    port map (
            O => \N__7348\,
            I => \N__7312\
        );

    \I__1661\ : LocalMux
    port map (
            O => \N__7345\,
            I => \N__7312\
        );

    \I__1660\ : Span4Mux_v
    port map (
            O => \N__7340\,
            I => \N__7305\
        );

    \I__1659\ : Span4Mux_v
    port map (
            O => \N__7329\,
            I => \N__7302\
        );

    \I__1658\ : InMux
    port map (
            O => \N__7328\,
            I => \N__7297\
        );

    \I__1657\ : InMux
    port map (
            O => \N__7327\,
            I => \N__7297\
        );

    \I__1656\ : InMux
    port map (
            O => \N__7324\,
            I => \N__7294\
        );

    \I__1655\ : Span12Mux_s2_v
    port map (
            O => \N__7321\,
            I => \N__7291\
        );

    \I__1654\ : Span4Mux_v
    port map (
            O => \N__7312\,
            I => \N__7288\
        );

    \I__1653\ : InMux
    port map (
            O => \N__7311\,
            I => \N__7285\
        );

    \I__1652\ : InMux
    port map (
            O => \N__7310\,
            I => \N__7278\
        );

    \I__1651\ : InMux
    port map (
            O => \N__7309\,
            I => \N__7278\
        );

    \I__1650\ : InMux
    port map (
            O => \N__7308\,
            I => \N__7278\
        );

    \I__1649\ : Sp12to4
    port map (
            O => \N__7305\,
            I => \N__7269\
        );

    \I__1648\ : Sp12to4
    port map (
            O => \N__7302\,
            I => \N__7269\
        );

    \I__1647\ : LocalMux
    port map (
            O => \N__7297\,
            I => \N__7269\
        );

    \I__1646\ : LocalMux
    port map (
            O => \N__7294\,
            I => \N__7269\
        );

    \I__1645\ : Odrv12
    port map (
            O => \N__7291\,
            I => \uut.inc\
        );

    \I__1644\ : Odrv4
    port map (
            O => \N__7288\,
            I => \uut.inc\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__7285\,
            I => \uut.inc\
        );

    \I__1642\ : LocalMux
    port map (
            O => \N__7278\,
            I => \uut.inc\
        );

    \I__1641\ : Odrv12
    port map (
            O => \N__7269\,
            I => \uut.inc\
        );

    \I__1640\ : CascadeMux
    port map (
            O => \N__7258\,
            I => \N__7255\
        );

    \I__1639\ : InMux
    port map (
            O => \N__7255\,
            I => \N__7251\
        );

    \I__1638\ : CascadeMux
    port map (
            O => \N__7254\,
            I => \N__7248\
        );

    \I__1637\ : LocalMux
    port map (
            O => \N__7251\,
            I => \N__7244\
        );

    \I__1636\ : InMux
    port map (
            O => \N__7248\,
            I => \N__7239\
        );

    \I__1635\ : InMux
    port map (
            O => \N__7247\,
            I => \N__7239\
        );

    \I__1634\ : Span4Mux_h
    port map (
            O => \N__7244\,
            I => \N__7234\
        );

    \I__1633\ : LocalMux
    port map (
            O => \N__7239\,
            I => \N__7231\
        );

    \I__1632\ : InMux
    port map (
            O => \N__7238\,
            I => \N__7228\
        );

    \I__1631\ : InMux
    port map (
            O => \N__7237\,
            I => \N__7225\
        );

    \I__1630\ : Span4Mux_v
    port map (
            O => \N__7234\,
            I => \N__7222\
        );

    \I__1629\ : Span12Mux_v
    port map (
            O => \N__7231\,
            I => \N__7217\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__7228\,
            I => \N__7217\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__7225\,
            I => \uut.ir_out_2\
        );

    \I__1626\ : Odrv4
    port map (
            O => \N__7222\,
            I => \uut.ir_out_2\
        );

    \I__1625\ : Odrv12
    port map (
            O => \N__7217\,
            I => \uut.ir_out_2\
        );

    \I__1624\ : InMux
    port map (
            O => \N__7210\,
            I => \N__7206\
        );

    \I__1623\ : InMux
    port map (
            O => \N__7209\,
            I => \N__7203\
        );

    \I__1622\ : LocalMux
    port map (
            O => \N__7206\,
            I => \N__7200\
        );

    \I__1621\ : LocalMux
    port map (
            O => \N__7203\,
            I => \N__7197\
        );

    \I__1620\ : Odrv4
    port map (
            O => \N__7200\,
            I => \uut.N_14_0\
        );

    \I__1619\ : Odrv4
    port map (
            O => \N__7197\,
            I => \uut.N_14_0\
        );

    \I__1618\ : InMux
    port map (
            O => \N__7192\,
            I => \N__7189\
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__7189\,
            I => \N__7186\
        );

    \I__1616\ : Span4Mux_s3_h
    port map (
            O => \N__7186\,
            I => \N__7182\
        );

    \I__1615\ : InMux
    port map (
            O => \N__7185\,
            I => \N__7179\
        );

    \I__1614\ : Odrv4
    port map (
            O => \N__7182\,
            I => \uut.alu_out_m_0_2\
        );

    \I__1613\ : LocalMux
    port map (
            O => \N__7179\,
            I => \uut.alu_out_m_0_2\
        );

    \I__1612\ : CascadeMux
    port map (
            O => \N__7174\,
            I => \uut.out_1_0_iv_3_cascade_\
        );

    \I__1611\ : CascadeMux
    port map (
            O => \N__7171\,
            I => \N__7168\
        );

    \I__1610\ : InMux
    port map (
            O => \N__7168\,
            I => \N__7164\
        );

    \I__1609\ : InMux
    port map (
            O => \N__7167\,
            I => \N__7160\
        );

    \I__1608\ : LocalMux
    port map (
            O => \N__7164\,
            I => \N__7157\
        );

    \I__1607\ : InMux
    port map (
            O => \N__7163\,
            I => \N__7154\
        );

    \I__1606\ : LocalMux
    port map (
            O => \N__7160\,
            I => \N__7151\
        );

    \I__1605\ : Span12Mux_s11_h
    port map (
            O => \N__7157\,
            I => \N__7148\
        );

    \I__1604\ : LocalMux
    port map (
            O => \N__7154\,
            I => \uut.AR_out_2\
        );

    \I__1603\ : Odrv12
    port map (
            O => \N__7151\,
            I => \uut.AR_out_2\
        );

    \I__1602\ : Odrv12
    port map (
            O => \N__7148\,
            I => \uut.AR_out_2\
        );

    \I__1601\ : InMux
    port map (
            O => \N__7141\,
            I => \N__7136\
        );

    \I__1600\ : InMux
    port map (
            O => \N__7140\,
            I => \N__7133\
        );

    \I__1599\ : InMux
    port map (
            O => \N__7139\,
            I => \N__7129\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__7136\,
            I => \N__7126\
        );

    \I__1597\ : LocalMux
    port map (
            O => \N__7133\,
            I => \N__7123\
        );

    \I__1596\ : InMux
    port map (
            O => \N__7132\,
            I => \N__7120\
        );

    \I__1595\ : LocalMux
    port map (
            O => \N__7129\,
            I => \N__7117\
        );

    \I__1594\ : Span4Mux_s2_h
    port map (
            O => \N__7126\,
            I => \N__7114\
        );

    \I__1593\ : Span4Mux_v
    port map (
            O => \N__7123\,
            I => \N__7109\
        );

    \I__1592\ : LocalMux
    port map (
            O => \N__7120\,
            I => \N__7109\
        );

    \I__1591\ : Odrv4
    port map (
            O => \N__7117\,
            I => \uut.un11_MAR_LD\
        );

    \I__1590\ : Odrv4
    port map (
            O => \N__7114\,
            I => \uut.un11_MAR_LD\
        );

    \I__1589\ : Odrv4
    port map (
            O => \N__7109\,
            I => \uut.un11_MAR_LD\
        );

    \I__1588\ : InMux
    port map (
            O => \N__7102\,
            I => \N__7099\
        );

    \I__1587\ : LocalMux
    port map (
            O => \N__7099\,
            I => \N__7096\
        );

    \I__1586\ : Span4Mux_h
    port map (
            O => \N__7096\,
            I => \N__7093\
        );

    \I__1585\ : Odrv4
    port map (
            O => \N__7093\,
            I => \uut.MAR_LD_1\
        );

    \I__1584\ : InMux
    port map (
            O => \N__7090\,
            I => \N__7087\
        );

    \I__1583\ : LocalMux
    port map (
            O => \N__7087\,
            I => \uut.seq.counter.MAR_LD_0_0\
        );

    \I__1582\ : CascadeMux
    port map (
            O => \N__7084\,
            I => \uut.MAR_LD_1_cascade_\
        );

    \I__1581\ : CascadeMux
    port map (
            O => \N__7081\,
            I => \N__7078\
        );

    \I__1580\ : InMux
    port map (
            O => \N__7078\,
            I => \N__7075\
        );

    \I__1579\ : LocalMux
    port map (
            O => \N__7075\,
            I => \uut.N_16_0\
        );

    \I__1578\ : InMux
    port map (
            O => \N__7072\,
            I => \N__7069\
        );

    \I__1577\ : LocalMux
    port map (
            O => \N__7069\,
            I => \N__7066\
        );

    \I__1576\ : Odrv4
    port map (
            O => \N__7066\,
            I => \uut.alu_out_m_1_3\
        );

    \I__1575\ : CascadeMux
    port map (
            O => \N__7063\,
            I => \uut.AR_BUF.g0Z0Z_5_cascade_\
        );

    \I__1574\ : InMux
    port map (
            O => \N__7060\,
            I => \N__7056\
        );

    \I__1573\ : CascadeMux
    port map (
            O => \N__7059\,
            I => \N__7053\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__7056\,
            I => \N__7050\
        );

    \I__1571\ : InMux
    port map (
            O => \N__7053\,
            I => \N__7046\
        );

    \I__1570\ : Span4Mux_s2_h
    port map (
            O => \N__7050\,
            I => \N__7043\
        );

    \I__1569\ : InMux
    port map (
            O => \N__7049\,
            I => \N__7040\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__7046\,
            I => \uut.seq.D_2_1\
        );

    \I__1567\ : Odrv4
    port map (
            O => \N__7043\,
            I => \uut.seq.D_2_1\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__7040\,
            I => \uut.seq.D_2_1\
        );

    \I__1565\ : InMux
    port map (
            O => \N__7033\,
            I => \N__7024\
        );

    \I__1564\ : InMux
    port map (
            O => \N__7032\,
            I => \N__7021\
        );

    \I__1563\ : CascadeMux
    port map (
            O => \N__7031\,
            I => \N__7016\
        );

    \I__1562\ : CascadeMux
    port map (
            O => \N__7030\,
            I => \N__7013\
        );

    \I__1561\ : InMux
    port map (
            O => \N__7029\,
            I => \N__7010\
        );

    \I__1560\ : InMux
    port map (
            O => \N__7028\,
            I => \N__7007\
        );

    \I__1559\ : InMux
    port map (
            O => \N__7027\,
            I => \N__7004\
        );

    \I__1558\ : LocalMux
    port map (
            O => \N__7024\,
            I => \N__7001\
        );

    \I__1557\ : LocalMux
    port map (
            O => \N__7021\,
            I => \N__6998\
        );

    \I__1556\ : InMux
    port map (
            O => \N__7020\,
            I => \N__6995\
        );

    \I__1555\ : InMux
    port map (
            O => \N__7019\,
            I => \N__6990\
        );

    \I__1554\ : InMux
    port map (
            O => \N__7016\,
            I => \N__6990\
        );

    \I__1553\ : InMux
    port map (
            O => \N__7013\,
            I => \N__6987\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__7010\,
            I => \N__6982\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__7007\,
            I => \N__6982\
        );

    \I__1550\ : LocalMux
    port map (
            O => \N__7004\,
            I => \N__6979\
        );

    \I__1549\ : Span4Mux_v
    port map (
            O => \N__7001\,
            I => \N__6976\
        );

    \I__1548\ : Span12Mux_s4_h
    port map (
            O => \N__6998\,
            I => \N__6971\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__6995\,
            I => \N__6971\
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__6990\,
            I => \N__6966\
        );

    \I__1545\ : LocalMux
    port map (
            O => \N__6987\,
            I => \N__6966\
        );

    \I__1544\ : Odrv4
    port map (
            O => \N__6982\,
            I => \uut.ir_out_i_2_6\
        );

    \I__1543\ : Odrv12
    port map (
            O => \N__6979\,
            I => \uut.ir_out_i_2_6\
        );

    \I__1542\ : Odrv4
    port map (
            O => \N__6976\,
            I => \uut.ir_out_i_2_6\
        );

    \I__1541\ : Odrv12
    port map (
            O => \N__6971\,
            I => \uut.ir_out_i_2_6\
        );

    \I__1540\ : Odrv4
    port map (
            O => \N__6966\,
            I => \uut.ir_out_i_2_6\
        );

    \I__1539\ : CascadeMux
    port map (
            O => \N__6955\,
            I => \N__6952\
        );

    \I__1538\ : InMux
    port map (
            O => \N__6952\,
            I => \N__6949\
        );

    \I__1537\ : LocalMux
    port map (
            O => \N__6949\,
            I => \N__6946\
        );

    \I__1536\ : Odrv4
    port map (
            O => \N__6946\,
            I => \uut.seq.D_2\
        );

    \I__1535\ : InMux
    port map (
            O => \N__6943\,
            I => \N__6939\
        );

    \I__1534\ : InMux
    port map (
            O => \N__6942\,
            I => \N__6936\
        );

    \I__1533\ : LocalMux
    port map (
            O => \N__6939\,
            I => \N__6931\
        );

    \I__1532\ : LocalMux
    port map (
            O => \N__6936\,
            I => \N__6928\
        );

    \I__1531\ : InMux
    port map (
            O => \N__6935\,
            I => \N__6922\
        );

    \I__1530\ : InMux
    port map (
            O => \N__6934\,
            I => \N__6919\
        );

    \I__1529\ : Span4Mux_s3_h
    port map (
            O => \N__6931\,
            I => \N__6916\
        );

    \I__1528\ : Span12Mux_s9_v
    port map (
            O => \N__6928\,
            I => \N__6913\
        );

    \I__1527\ : InMux
    port map (
            O => \N__6927\,
            I => \N__6908\
        );

    \I__1526\ : InMux
    port map (
            O => \N__6926\,
            I => \N__6908\
        );

    \I__1525\ : InMux
    port map (
            O => \N__6925\,
            I => \N__6905\
        );

    \I__1524\ : LocalMux
    port map (
            O => \N__6922\,
            I => \uut.ir_out_i_2_5\
        );

    \I__1523\ : LocalMux
    port map (
            O => \N__6919\,
            I => \uut.ir_out_i_2_5\
        );

    \I__1522\ : Odrv4
    port map (
            O => \N__6916\,
            I => \uut.ir_out_i_2_5\
        );

    \I__1521\ : Odrv12
    port map (
            O => \N__6913\,
            I => \uut.ir_out_i_2_5\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__6908\,
            I => \uut.ir_out_i_2_5\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__6905\,
            I => \uut.ir_out_i_2_5\
        );

    \I__1518\ : CascadeMux
    port map (
            O => \N__6892\,
            I => \uut.B_LD_0_1_tz_cascade_\
        );

    \I__1517\ : InMux
    port map (
            O => \N__6889\,
            I => \N__6886\
        );

    \I__1516\ : LocalMux
    port map (
            O => \N__6886\,
            I => \N__6881\
        );

    \I__1515\ : InMux
    port map (
            O => \N__6885\,
            I => \N__6878\
        );

    \I__1514\ : CascadeMux
    port map (
            O => \N__6884\,
            I => \N__6875\
        );

    \I__1513\ : Span4Mux_h
    port map (
            O => \N__6881\,
            I => \N__6869\
        );

    \I__1512\ : LocalMux
    port map (
            O => \N__6878\,
            I => \N__6869\
        );

    \I__1511\ : InMux
    port map (
            O => \N__6875\,
            I => \N__6866\
        );

    \I__1510\ : InMux
    port map (
            O => \N__6874\,
            I => \N__6863\
        );

    \I__1509\ : Span4Mux_h
    port map (
            O => \N__6869\,
            I => \N__6860\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__6866\,
            I => \N__6857\
        );

    \I__1507\ : LocalMux
    port map (
            O => \N__6863\,
            I => \N__6854\
        );

    \I__1506\ : Odrv4
    port map (
            O => \N__6860\,
            I => \uut.mem.i2_mux_0\
        );

    \I__1505\ : Odrv12
    port map (
            O => \N__6857\,
            I => \uut.mem.i2_mux_0\
        );

    \I__1504\ : Odrv12
    port map (
            O => \N__6854\,
            I => \uut.mem.i2_mux_0\
        );

    \I__1503\ : InMux
    port map (
            O => \N__6847\,
            I => \N__6844\
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__6844\,
            I => \N__6841\
        );

    \I__1501\ : Odrv12
    port map (
            O => \N__6841\,
            I => \uut.out_1_0_iv_2_1\
        );

    \I__1500\ : IoInMux
    port map (
            O => \N__6838\,
            I => \N__6835\
        );

    \I__1499\ : LocalMux
    port map (
            O => \N__6835\,
            I => \N__6831\
        );

    \I__1498\ : CascadeMux
    port map (
            O => \N__6834\,
            I => \N__6828\
        );

    \I__1497\ : IoSpan4Mux
    port map (
            O => \N__6831\,
            I => \N__6825\
        );

    \I__1496\ : InMux
    port map (
            O => \N__6828\,
            I => \N__6822\
        );

    \I__1495\ : Odrv4
    port map (
            O => \N__6825\,
            I => \LED3_c\
        );

    \I__1494\ : LocalMux
    port map (
            O => \N__6822\,
            I => \LED3_c\
        );

    \I__1493\ : InMux
    port map (
            O => \N__6817\,
            I => \N__6814\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__6814\,
            I => \N__6811\
        );

    \I__1491\ : Span4Mux_h
    port map (
            O => \N__6811\,
            I => \N__6808\
        );

    \I__1490\ : Span4Mux_v
    port map (
            O => \N__6808\,
            I => \N__6805\
        );

    \I__1489\ : Odrv4
    port map (
            O => \N__6805\,
            I => \uut.m10\
        );

    \I__1488\ : CascadeMux
    port map (
            O => \N__6802\,
            I => \uut.m10_cascade_\
        );

    \I__1487\ : InMux
    port map (
            O => \N__6799\,
            I => \N__6795\
        );

    \I__1486\ : InMux
    port map (
            O => \N__6798\,
            I => \N__6792\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__6795\,
            I => \N__6789\
        );

    \I__1484\ : LocalMux
    port map (
            O => \N__6792\,
            I => \N__6786\
        );

    \I__1483\ : Span4Mux_s1_v
    port map (
            O => \N__6789\,
            I => \N__6783\
        );

    \I__1482\ : Span4Mux_h
    port map (
            O => \N__6786\,
            I => \N__6780\
        );

    \I__1481\ : Odrv4
    port map (
            O => \N__6783\,
            I => \uut.b_reg_out_0\
        );

    \I__1480\ : Odrv4
    port map (
            O => \N__6780\,
            I => \uut.b_reg_out_0\
        );

    \I__1479\ : InMux
    port map (
            O => \N__6775\,
            I => \N__6769\
        );

    \I__1478\ : InMux
    port map (
            O => \N__6774\,
            I => \N__6763\
        );

    \I__1477\ : InMux
    port map (
            O => \N__6773\,
            I => \N__6755\
        );

    \I__1476\ : InMux
    port map (
            O => \N__6772\,
            I => \N__6755\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__6769\,
            I => \N__6749\
        );

    \I__1474\ : InMux
    port map (
            O => \N__6768\,
            I => \N__6746\
        );

    \I__1473\ : InMux
    port map (
            O => \N__6767\,
            I => \N__6743\
        );

    \I__1472\ : InMux
    port map (
            O => \N__6766\,
            I => \N__6740\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__6763\,
            I => \N__6737\
        );

    \I__1470\ : InMux
    port map (
            O => \N__6762\,
            I => \N__6732\
        );

    \I__1469\ : InMux
    port map (
            O => \N__6761\,
            I => \N__6732\
        );

    \I__1468\ : InMux
    port map (
            O => \N__6760\,
            I => \N__6729\
        );

    \I__1467\ : LocalMux
    port map (
            O => \N__6755\,
            I => \N__6726\
        );

    \I__1466\ : InMux
    port map (
            O => \N__6754\,
            I => \N__6723\
        );

    \I__1465\ : InMux
    port map (
            O => \N__6753\,
            I => \N__6718\
        );

    \I__1464\ : InMux
    port map (
            O => \N__6752\,
            I => \N__6718\
        );

    \I__1463\ : Span4Mux_v
    port map (
            O => \N__6749\,
            I => \N__6713\
        );

    \I__1462\ : LocalMux
    port map (
            O => \N__6746\,
            I => \N__6713\
        );

    \I__1461\ : LocalMux
    port map (
            O => \N__6743\,
            I => \N__6706\
        );

    \I__1460\ : LocalMux
    port map (
            O => \N__6740\,
            I => \N__6706\
        );

    \I__1459\ : Span4Mux_v
    port map (
            O => \N__6737\,
            I => \N__6706\
        );

    \I__1458\ : LocalMux
    port map (
            O => \N__6732\,
            I => \N__6703\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__6729\,
            I => \N__6700\
        );

    \I__1456\ : Span4Mux_s3_h
    port map (
            O => \N__6726\,
            I => \N__6693\
        );

    \I__1455\ : LocalMux
    port map (
            O => \N__6723\,
            I => \N__6693\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__6718\,
            I => \N__6693\
        );

    \I__1453\ : Span4Mux_v
    port map (
            O => \N__6713\,
            I => \N__6690\
        );

    \I__1452\ : Span4Mux_h
    port map (
            O => \N__6706\,
            I => \N__6685\
        );

    \I__1451\ : Span4Mux_s2_h
    port map (
            O => \N__6703\,
            I => \N__6685\
        );

    \I__1450\ : Span4Mux_h
    port map (
            O => \N__6700\,
            I => \N__6680\
        );

    \I__1449\ : Span4Mux_v
    port map (
            O => \N__6693\,
            I => \N__6680\
        );

    \I__1448\ : Odrv4
    port map (
            O => \N__6690\,
            I => \uut.T_1_fast_RNI28LI1_0\
        );

    \I__1447\ : Odrv4
    port map (
            O => \N__6685\,
            I => \uut.T_1_fast_RNI28LI1_0\
        );

    \I__1446\ : Odrv4
    port map (
            O => \N__6680\,
            I => \uut.T_1_fast_RNI28LI1_0\
        );

    \I__1445\ : CascadeMux
    port map (
            O => \N__6673\,
            I => \N__6669\
        );

    \I__1444\ : InMux
    port map (
            O => \N__6672\,
            I => \N__6665\
        );

    \I__1443\ : InMux
    port map (
            O => \N__6669\,
            I => \N__6660\
        );

    \I__1442\ : InMux
    port map (
            O => \N__6668\,
            I => \N__6660\
        );

    \I__1441\ : LocalMux
    port map (
            O => \N__6665\,
            I => \N__6657\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__6660\,
            I => \N__6654\
        );

    \I__1439\ : Span4Mux_s2_h
    port map (
            O => \N__6657\,
            I => \N__6650\
        );

    \I__1438\ : Span4Mux_s2_h
    port map (
            O => \N__6654\,
            I => \N__6647\
        );

    \I__1437\ : InMux
    port map (
            O => \N__6653\,
            I => \N__6644\
        );

    \I__1436\ : Odrv4
    port map (
            O => \N__6650\,
            I => \uut.b_reg_out_3\
        );

    \I__1435\ : Odrv4
    port map (
            O => \N__6647\,
            I => \uut.b_reg_out_3\
        );

    \I__1434\ : LocalMux
    port map (
            O => \N__6644\,
            I => \uut.b_reg_out_3\
        );

    \I__1433\ : InMux
    port map (
            O => \N__6637\,
            I => \N__6628\
        );

    \I__1432\ : InMux
    port map (
            O => \N__6636\,
            I => \N__6628\
        );

    \I__1431\ : InMux
    port map (
            O => \N__6635\,
            I => \N__6628\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__6628\,
            I => \N__6625\
        );

    \I__1429\ : Odrv4
    port map (
            O => \N__6625\,
            I => \uut.un1_A_cry_2_c_RNIBSP45\
        );

    \I__1428\ : InMux
    port map (
            O => \N__6622\,
            I => \N__6611\
        );

    \I__1427\ : InMux
    port map (
            O => \N__6621\,
            I => \N__6607\
        );

    \I__1426\ : InMux
    port map (
            O => \N__6620\,
            I => \N__6604\
        );

    \I__1425\ : InMux
    port map (
            O => \N__6619\,
            I => \N__6600\
        );

    \I__1424\ : InMux
    port map (
            O => \N__6618\,
            I => \N__6597\
        );

    \I__1423\ : InMux
    port map (
            O => \N__6617\,
            I => \N__6594\
        );

    \I__1422\ : InMux
    port map (
            O => \N__6616\,
            I => \N__6591\
        );

    \I__1421\ : InMux
    port map (
            O => \N__6615\,
            I => \N__6586\
        );

    \I__1420\ : InMux
    port map (
            O => \N__6614\,
            I => \N__6586\
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__6611\,
            I => \N__6583\
        );

    \I__1418\ : CascadeMux
    port map (
            O => \N__6610\,
            I => \N__6577\
        );

    \I__1417\ : LocalMux
    port map (
            O => \N__6607\,
            I => \N__6572\
        );

    \I__1416\ : LocalMux
    port map (
            O => \N__6604\,
            I => \N__6572\
        );

    \I__1415\ : CascadeMux
    port map (
            O => \N__6603\,
            I => \N__6569\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__6600\,
            I => \N__6566\
        );

    \I__1413\ : LocalMux
    port map (
            O => \N__6597\,
            I => \N__6563\
        );

    \I__1412\ : LocalMux
    port map (
            O => \N__6594\,
            I => \N__6560\
        );

    \I__1411\ : LocalMux
    port map (
            O => \N__6591\,
            I => \N__6557\
        );

    \I__1410\ : LocalMux
    port map (
            O => \N__6586\,
            I => \N__6554\
        );

    \I__1409\ : Span4Mux_v
    port map (
            O => \N__6583\,
            I => \N__6551\
        );

    \I__1408\ : InMux
    port map (
            O => \N__6582\,
            I => \N__6548\
        );

    \I__1407\ : InMux
    port map (
            O => \N__6581\,
            I => \N__6543\
        );

    \I__1406\ : InMux
    port map (
            O => \N__6580\,
            I => \N__6543\
        );

    \I__1405\ : InMux
    port map (
            O => \N__6577\,
            I => \N__6540\
        );

    \I__1404\ : Span4Mux_h
    port map (
            O => \N__6572\,
            I => \N__6537\
        );

    \I__1403\ : InMux
    port map (
            O => \N__6569\,
            I => \N__6534\
        );

    \I__1402\ : Span4Mux_h
    port map (
            O => \N__6566\,
            I => \N__6531\
        );

    \I__1401\ : Span4Mux_v
    port map (
            O => \N__6563\,
            I => \N__6516\
        );

    \I__1400\ : Span4Mux_v
    port map (
            O => \N__6560\,
            I => \N__6516\
        );

    \I__1399\ : Span4Mux_h
    port map (
            O => \N__6557\,
            I => \N__6516\
        );

    \I__1398\ : Span4Mux_v
    port map (
            O => \N__6554\,
            I => \N__6516\
        );

    \I__1397\ : Span4Mux_s0_h
    port map (
            O => \N__6551\,
            I => \N__6516\
        );

    \I__1396\ : LocalMux
    port map (
            O => \N__6548\,
            I => \N__6516\
        );

    \I__1395\ : LocalMux
    port map (
            O => \N__6543\,
            I => \N__6516\
        );

    \I__1394\ : LocalMux
    port map (
            O => \N__6540\,
            I => \uut.un1_ALU_en_0\
        );

    \I__1393\ : Odrv4
    port map (
            O => \N__6537\,
            I => \uut.un1_ALU_en_0\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__6534\,
            I => \uut.un1_ALU_en_0\
        );

    \I__1391\ : Odrv4
    port map (
            O => \N__6531\,
            I => \uut.un1_ALU_en_0\
        );

    \I__1390\ : Odrv4
    port map (
            O => \N__6516\,
            I => \uut.un1_ALU_en_0\
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__6505\,
            I => \uut.ALU_main.N_44_cascade_\
        );

    \I__1388\ : InMux
    port map (
            O => \N__6502\,
            I => \N__6493\
        );

    \I__1387\ : InMux
    port map (
            O => \N__6501\,
            I => \N__6489\
        );

    \I__1386\ : InMux
    port map (
            O => \N__6500\,
            I => \N__6486\
        );

    \I__1385\ : InMux
    port map (
            O => \N__6499\,
            I => \N__6479\
        );

    \I__1384\ : InMux
    port map (
            O => \N__6498\,
            I => \N__6479\
        );

    \I__1383\ : InMux
    port map (
            O => \N__6497\,
            I => \N__6479\
        );

    \I__1382\ : CascadeMux
    port map (
            O => \N__6496\,
            I => \N__6476\
        );

    \I__1381\ : LocalMux
    port map (
            O => \N__6493\,
            I => \N__6471\
        );

    \I__1380\ : InMux
    port map (
            O => \N__6492\,
            I => \N__6468\
        );

    \I__1379\ : LocalMux
    port map (
            O => \N__6489\,
            I => \N__6464\
        );

    \I__1378\ : LocalMux
    port map (
            O => \N__6486\,
            I => \N__6460\
        );

    \I__1377\ : LocalMux
    port map (
            O => \N__6479\,
            I => \N__6457\
        );

    \I__1376\ : InMux
    port map (
            O => \N__6476\,
            I => \N__6453\
        );

    \I__1375\ : InMux
    port map (
            O => \N__6475\,
            I => \N__6450\
        );

    \I__1374\ : InMux
    port map (
            O => \N__6474\,
            I => \N__6447\
        );

    \I__1373\ : Span4Mux_v
    port map (
            O => \N__6471\,
            I => \N__6442\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__6468\,
            I => \N__6442\
        );

    \I__1371\ : InMux
    port map (
            O => \N__6467\,
            I => \N__6439\
        );

    \I__1370\ : Span4Mux_h
    port map (
            O => \N__6464\,
            I => \N__6436\
        );

    \I__1369\ : InMux
    port map (
            O => \N__6463\,
            I => \N__6433\
        );

    \I__1368\ : Span4Mux_v
    port map (
            O => \N__6460\,
            I => \N__6428\
        );

    \I__1367\ : Span4Mux_v
    port map (
            O => \N__6457\,
            I => \N__6428\
        );

    \I__1366\ : InMux
    port map (
            O => \N__6456\,
            I => \N__6425\
        );

    \I__1365\ : LocalMux
    port map (
            O => \N__6453\,
            I => \uut.T_1_fast_RNIVM0N3_0\
        );

    \I__1364\ : LocalMux
    port map (
            O => \N__6450\,
            I => \uut.T_1_fast_RNIVM0N3_0\
        );

    \I__1363\ : LocalMux
    port map (
            O => \N__6447\,
            I => \uut.T_1_fast_RNIVM0N3_0\
        );

    \I__1362\ : Odrv4
    port map (
            O => \N__6442\,
            I => \uut.T_1_fast_RNIVM0N3_0\
        );

    \I__1361\ : LocalMux
    port map (
            O => \N__6439\,
            I => \uut.T_1_fast_RNIVM0N3_0\
        );

    \I__1360\ : Odrv4
    port map (
            O => \N__6436\,
            I => \uut.T_1_fast_RNIVM0N3_0\
        );

    \I__1359\ : LocalMux
    port map (
            O => \N__6433\,
            I => \uut.T_1_fast_RNIVM0N3_0\
        );

    \I__1358\ : Odrv4
    port map (
            O => \N__6428\,
            I => \uut.T_1_fast_RNIVM0N3_0\
        );

    \I__1357\ : LocalMux
    port map (
            O => \N__6425\,
            I => \uut.T_1_fast_RNIVM0N3_0\
        );

    \I__1356\ : InMux
    port map (
            O => \N__6406\,
            I => \N__6403\
        );

    \I__1355\ : LocalMux
    port map (
            O => \N__6403\,
            I => \N__6399\
        );

    \I__1354\ : InMux
    port map (
            O => \N__6402\,
            I => \N__6396\
        );

    \I__1353\ : Span4Mux_s1_h
    port map (
            O => \N__6399\,
            I => \N__6392\
        );

    \I__1352\ : LocalMux
    port map (
            O => \N__6396\,
            I => \N__6389\
        );

    \I__1351\ : InMux
    port map (
            O => \N__6395\,
            I => \N__6385\
        );

    \I__1350\ : Span4Mux_h
    port map (
            O => \N__6392\,
            I => \N__6380\
        );

    \I__1349\ : Span4Mux_h
    port map (
            O => \N__6389\,
            I => \N__6380\
        );

    \I__1348\ : InMux
    port map (
            O => \N__6388\,
            I => \N__6377\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__6385\,
            I => \N__6374\
        );

    \I__1346\ : Odrv4
    port map (
            O => \N__6380\,
            I => \uut.acc_out_m_6\
        );

    \I__1345\ : LocalMux
    port map (
            O => \N__6377\,
            I => \uut.acc_out_m_6\
        );

    \I__1344\ : Odrv12
    port map (
            O => \N__6374\,
            I => \uut.acc_out_m_6\
        );

    \I__1343\ : InMux
    port map (
            O => \N__6367\,
            I => \N__6364\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__6364\,
            I => \N__6360\
        );

    \I__1341\ : InMux
    port map (
            O => \N__6363\,
            I => \N__6356\
        );

    \I__1340\ : Span4Mux_v
    port map (
            O => \N__6360\,
            I => \N__6353\
        );

    \I__1339\ : InMux
    port map (
            O => \N__6359\,
            I => \N__6350\
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__6356\,
            I => \N__6346\
        );

    \I__1337\ : Span4Mux_h
    port map (
            O => \N__6353\,
            I => \N__6341\
        );

    \I__1336\ : LocalMux
    port map (
            O => \N__6350\,
            I => \N__6341\
        );

    \I__1335\ : InMux
    port map (
            O => \N__6349\,
            I => \N__6338\
        );

    \I__1334\ : Odrv4
    port map (
            O => \N__6346\,
            I => \uut.alu_out_m_6\
        );

    \I__1333\ : Odrv4
    port map (
            O => \N__6341\,
            I => \uut.alu_out_m_6\
        );

    \I__1332\ : LocalMux
    port map (
            O => \N__6338\,
            I => \uut.alu_out_m_6\
        );

    \I__1331\ : CascadeMux
    port map (
            O => \N__6331\,
            I => \N__6327\
        );

    \I__1330\ : CascadeMux
    port map (
            O => \N__6330\,
            I => \N__6324\
        );

    \I__1329\ : InMux
    port map (
            O => \N__6327\,
            I => \N__6321\
        );

    \I__1328\ : InMux
    port map (
            O => \N__6324\,
            I => \N__6317\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__6321\,
            I => \N__6313\
        );

    \I__1326\ : CascadeMux
    port map (
            O => \N__6320\,
            I => \N__6310\
        );

    \I__1325\ : LocalMux
    port map (
            O => \N__6317\,
            I => \N__6307\
        );

    \I__1324\ : CascadeMux
    port map (
            O => \N__6316\,
            I => \N__6304\
        );

    \I__1323\ : Span4Mux_v
    port map (
            O => \N__6313\,
            I => \N__6301\
        );

    \I__1322\ : InMux
    port map (
            O => \N__6310\,
            I => \N__6298\
        );

    \I__1321\ : Span4Mux_v
    port map (
            O => \N__6307\,
            I => \N__6295\
        );

    \I__1320\ : InMux
    port map (
            O => \N__6304\,
            I => \N__6292\
        );

    \I__1319\ : Span4Mux_h
    port map (
            O => \N__6301\,
            I => \N__6289\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__6298\,
            I => \N__6286\
        );

    \I__1317\ : Sp12to4
    port map (
            O => \N__6295\,
            I => \N__6281\
        );

    \I__1316\ : LocalMux
    port map (
            O => \N__6292\,
            I => \N__6281\
        );

    \I__1315\ : Odrv4
    port map (
            O => \N__6289\,
            I => \uut.mem.N_29_mux\
        );

    \I__1314\ : Odrv4
    port map (
            O => \N__6286\,
            I => \uut.mem.N_29_mux\
        );

    \I__1313\ : Odrv12
    port map (
            O => \N__6281\,
            I => \uut.mem.N_29_mux\
        );

    \I__1312\ : CascadeMux
    port map (
            O => \N__6274\,
            I => \N__6269\
        );

    \I__1311\ : InMux
    port map (
            O => \N__6273\,
            I => \N__6266\
        );

    \I__1310\ : InMux
    port map (
            O => \N__6272\,
            I => \N__6262\
        );

    \I__1309\ : InMux
    port map (
            O => \N__6269\,
            I => \N__6259\
        );

    \I__1308\ : LocalMux
    port map (
            O => \N__6266\,
            I => \N__6256\
        );

    \I__1307\ : InMux
    port map (
            O => \N__6265\,
            I => \N__6253\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__6262\,
            I => \N__6250\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__6259\,
            I => \N__6247\
        );

    \I__1304\ : Span4Mux_h
    port map (
            O => \N__6256\,
            I => \N__6244\
        );

    \I__1303\ : LocalMux
    port map (
            O => \N__6253\,
            I => \N__6239\
        );

    \I__1302\ : Span12Mux_v
    port map (
            O => \N__6250\,
            I => \N__6239\
        );

    \I__1301\ : Span4Mux_v
    port map (
            O => \N__6247\,
            I => \N__6236\
        );

    \I__1300\ : Odrv4
    port map (
            O => \N__6244\,
            I => \uut.acc_out_6\
        );

    \I__1299\ : Odrv12
    port map (
            O => \N__6239\,
            I => \uut.acc_out_6\
        );

    \I__1298\ : Odrv4
    port map (
            O => \N__6236\,
            I => \uut.acc_out_6\
        );

    \I__1297\ : CascadeMux
    port map (
            O => \N__6229\,
            I => \N__6225\
        );

    \I__1296\ : InMux
    port map (
            O => \N__6228\,
            I => \N__6222\
        );

    \I__1295\ : InMux
    port map (
            O => \N__6225\,
            I => \N__6219\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__6222\,
            I => \N__6216\
        );

    \I__1293\ : LocalMux
    port map (
            O => \N__6219\,
            I => \N__6210\
        );

    \I__1292\ : Span4Mux_s1_h
    port map (
            O => \N__6216\,
            I => \N__6210\
        );

    \I__1291\ : InMux
    port map (
            O => \N__6215\,
            I => \N__6207\
        );

    \I__1290\ : Span4Mux_h
    port map (
            O => \N__6210\,
            I => \N__6204\
        );

    \I__1289\ : LocalMux
    port map (
            O => \N__6207\,
            I => \uut.acc_out_m_7\
        );

    \I__1288\ : Odrv4
    port map (
            O => \N__6204\,
            I => \uut.acc_out_m_7\
        );

    \I__1287\ : InMux
    port map (
            O => \N__6199\,
            I => \N__6196\
        );

    \I__1286\ : LocalMux
    port map (
            O => \N__6196\,
            I => \N__6191\
        );

    \I__1285\ : InMux
    port map (
            O => \N__6195\,
            I => \N__6188\
        );

    \I__1284\ : InMux
    port map (
            O => \N__6194\,
            I => \N__6185\
        );

    \I__1283\ : Odrv12
    port map (
            O => \N__6191\,
            I => \uut.alu_out_m_7\
        );

    \I__1282\ : LocalMux
    port map (
            O => \N__6188\,
            I => \uut.alu_out_m_7\
        );

    \I__1281\ : LocalMux
    port map (
            O => \N__6185\,
            I => \uut.alu_out_m_7\
        );

    \I__1280\ : InMux
    port map (
            O => \N__6178\,
            I => \N__6174\
        );

    \I__1279\ : InMux
    port map (
            O => \N__6177\,
            I => \N__6171\
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__6174\,
            I => \N__6165\
        );

    \I__1277\ : LocalMux
    port map (
            O => \N__6171\,
            I => \N__6165\
        );

    \I__1276\ : InMux
    port map (
            O => \N__6170\,
            I => \N__6162\
        );

    \I__1275\ : Span4Mux_s3_v
    port map (
            O => \N__6165\,
            I => \N__6159\
        );

    \I__1274\ : LocalMux
    port map (
            O => \N__6162\,
            I => \N__6156\
        );

    \I__1273\ : Span4Mux_h
    port map (
            O => \N__6159\,
            I => \N__6153\
        );

    \I__1272\ : Span4Mux_h
    port map (
            O => \N__6156\,
            I => \N__6150\
        );

    \I__1271\ : Odrv4
    port map (
            O => \N__6153\,
            I => \uut.acc_out_7\
        );

    \I__1270\ : Odrv4
    port map (
            O => \N__6150\,
            I => \uut.acc_out_7\
        );

    \I__1269\ : InMux
    port map (
            O => \N__6145\,
            I => \N__6142\
        );

    \I__1268\ : LocalMux
    port map (
            O => \N__6142\,
            I => \N__6138\
        );

    \I__1267\ : InMux
    port map (
            O => \N__6141\,
            I => \N__6135\
        );

    \I__1266\ : Span4Mux_v
    port map (
            O => \N__6138\,
            I => \N__6132\
        );

    \I__1265\ : LocalMux
    port map (
            O => \N__6135\,
            I => \N__6129\
        );

    \I__1264\ : Span4Mux_h
    port map (
            O => \N__6132\,
            I => \N__6123\
        );

    \I__1263\ : Span4Mux_v
    port map (
            O => \N__6129\,
            I => \N__6123\
        );

    \I__1262\ : InMux
    port map (
            O => \N__6128\,
            I => \N__6120\
        );

    \I__1261\ : Odrv4
    port map (
            O => \N__6123\,
            I => \uut.alu_out_m_5\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__6120\,
            I => \uut.alu_out_m_5\
        );

    \I__1259\ : InMux
    port map (
            O => \N__6115\,
            I => \N__6111\
        );

    \I__1258\ : InMux
    port map (
            O => \N__6114\,
            I => \N__6108\
        );

    \I__1257\ : LocalMux
    port map (
            O => \N__6111\,
            I => \N__6105\
        );

    \I__1256\ : LocalMux
    port map (
            O => \N__6108\,
            I => \N__6102\
        );

    \I__1255\ : Span12Mux_s6_h
    port map (
            O => \N__6105\,
            I => \N__6097\
        );

    \I__1254\ : Span4Mux_v
    port map (
            O => \N__6102\,
            I => \N__6094\
        );

    \I__1253\ : InMux
    port map (
            O => \N__6101\,
            I => \N__6091\
        );

    \I__1252\ : InMux
    port map (
            O => \N__6100\,
            I => \N__6088\
        );

    \I__1251\ : Odrv12
    port map (
            O => \N__6097\,
            I => \uut.acc_out_m_5\
        );

    \I__1250\ : Odrv4
    port map (
            O => \N__6094\,
            I => \uut.acc_out_m_5\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__6091\,
            I => \uut.acc_out_m_5\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__6088\,
            I => \uut.acc_out_m_5\
        );

    \I__1247\ : CascadeMux
    port map (
            O => \N__6079\,
            I => \N__6075\
        );

    \I__1246\ : InMux
    port map (
            O => \N__6078\,
            I => \N__6071\
        );

    \I__1245\ : InMux
    port map (
            O => \N__6075\,
            I => \N__6067\
        );

    \I__1244\ : InMux
    port map (
            O => \N__6074\,
            I => \N__6064\
        );

    \I__1243\ : LocalMux
    port map (
            O => \N__6071\,
            I => \N__6061\
        );

    \I__1242\ : CascadeMux
    port map (
            O => \N__6070\,
            I => \N__6058\
        );

    \I__1241\ : LocalMux
    port map (
            O => \N__6067\,
            I => \N__6053\
        );

    \I__1240\ : LocalMux
    port map (
            O => \N__6064\,
            I => \N__6053\
        );

    \I__1239\ : Span4Mux_h
    port map (
            O => \N__6061\,
            I => \N__6050\
        );

    \I__1238\ : InMux
    port map (
            O => \N__6058\,
            I => \N__6047\
        );

    \I__1237\ : Span4Mux_h
    port map (
            O => \N__6053\,
            I => \N__6044\
        );

    \I__1236\ : Sp12to4
    port map (
            O => \N__6050\,
            I => \N__6039\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__6047\,
            I => \N__6039\
        );

    \I__1234\ : Span4Mux_h
    port map (
            O => \N__6044\,
            I => \N__6036\
        );

    \I__1233\ : Odrv12
    port map (
            O => \N__6039\,
            I => \uut.mem.m20\
        );

    \I__1232\ : Odrv4
    port map (
            O => \N__6036\,
            I => \uut.mem.m20\
        );

    \I__1231\ : CascadeMux
    port map (
            O => \N__6031\,
            I => \N__6025\
        );

    \I__1230\ : InMux
    port map (
            O => \N__6030\,
            I => \N__6022\
        );

    \I__1229\ : InMux
    port map (
            O => \N__6029\,
            I => \N__6019\
        );

    \I__1228\ : CascadeMux
    port map (
            O => \N__6028\,
            I => \N__6016\
        );

    \I__1227\ : InMux
    port map (
            O => \N__6025\,
            I => \N__6013\
        );

    \I__1226\ : LocalMux
    port map (
            O => \N__6022\,
            I => \N__6010\
        );

    \I__1225\ : LocalMux
    port map (
            O => \N__6019\,
            I => \N__6007\
        );

    \I__1224\ : InMux
    port map (
            O => \N__6016\,
            I => \N__6004\
        );

    \I__1223\ : LocalMux
    port map (
            O => \N__6013\,
            I => \N__6001\
        );

    \I__1222\ : Span4Mux_v
    port map (
            O => \N__6010\,
            I => \N__5994\
        );

    \I__1221\ : Span4Mux_h
    port map (
            O => \N__6007\,
            I => \N__5994\
        );

    \I__1220\ : LocalMux
    port map (
            O => \N__6004\,
            I => \N__5994\
        );

    \I__1219\ : Span4Mux_h
    port map (
            O => \N__6001\,
            I => \N__5991\
        );

    \I__1218\ : Span4Mux_h
    port map (
            O => \N__5994\,
            I => \N__5988\
        );

    \I__1217\ : Odrv4
    port map (
            O => \N__5991\,
            I => \uut.acc_out_5\
        );

    \I__1216\ : Odrv4
    port map (
            O => \N__5988\,
            I => \uut.acc_out_5\
        );

    \I__1215\ : CascadeMux
    port map (
            O => \N__5983\,
            I => \N__5980\
        );

    \I__1214\ : InMux
    port map (
            O => \N__5980\,
            I => \N__5976\
        );

    \I__1213\ : InMux
    port map (
            O => \N__5979\,
            I => \N__5973\
        );

    \I__1212\ : LocalMux
    port map (
            O => \N__5976\,
            I => \N__5970\
        );

    \I__1211\ : LocalMux
    port map (
            O => \N__5973\,
            I => \N__5967\
        );

    \I__1210\ : Span4Mux_v
    port map (
            O => \N__5970\,
            I => \N__5961\
        );

    \I__1209\ : Span4Mux_v
    port map (
            O => \N__5967\,
            I => \N__5961\
        );

    \I__1208\ : InMux
    port map (
            O => \N__5966\,
            I => \N__5958\
        );

    \I__1207\ : Odrv4
    port map (
            O => \N__5961\,
            I => \uut.q_RNIDGA71\
        );

    \I__1206\ : LocalMux
    port map (
            O => \N__5958\,
            I => \uut.q_RNIDGA71\
        );

    \I__1205\ : CascadeMux
    port map (
            O => \N__5953\,
            I => \N__5950\
        );

    \I__1204\ : InMux
    port map (
            O => \N__5950\,
            I => \N__5943\
        );

    \I__1203\ : InMux
    port map (
            O => \N__5949\,
            I => \N__5940\
        );

    \I__1202\ : InMux
    port map (
            O => \N__5948\,
            I => \N__5933\
        );

    \I__1201\ : InMux
    port map (
            O => \N__5947\,
            I => \N__5933\
        );

    \I__1200\ : InMux
    port map (
            O => \N__5946\,
            I => \N__5933\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__5943\,
            I => \N__5930\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__5940\,
            I => \N__5925\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__5933\,
            I => \N__5925\
        );

    \I__1196\ : Span4Mux_v
    port map (
            O => \N__5930\,
            I => \N__5920\
        );

    \I__1195\ : Span4Mux_v
    port map (
            O => \N__5925\,
            I => \N__5920\
        );

    \I__1194\ : Odrv4
    port map (
            O => \N__5920\,
            I => \uut.mem.i2_mux\
        );

    \I__1193\ : InMux
    port map (
            O => \N__5917\,
            I => \N__5914\
        );

    \I__1192\ : LocalMux
    port map (
            O => \N__5914\,
            I => \N__5910\
        );

    \I__1191\ : InMux
    port map (
            O => \N__5913\,
            I => \N__5907\
        );

    \I__1190\ : Span4Mux_v
    port map (
            O => \N__5910\,
            I => \N__5902\
        );

    \I__1189\ : LocalMux
    port map (
            O => \N__5907\,
            I => \N__5899\
        );

    \I__1188\ : InMux
    port map (
            O => \N__5906\,
            I => \N__5896\
        );

    \I__1187\ : InMux
    port map (
            O => \N__5905\,
            I => \N__5893\
        );

    \I__1186\ : Odrv4
    port map (
            O => \N__5902\,
            I => \uut.alu_out_m_4\
        );

    \I__1185\ : Odrv4
    port map (
            O => \N__5899\,
            I => \uut.alu_out_m_4\
        );

    \I__1184\ : LocalMux
    port map (
            O => \N__5896\,
            I => \uut.alu_out_m_4\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__5893\,
            I => \uut.alu_out_m_4\
        );

    \I__1182\ : CascadeMux
    port map (
            O => \N__5884\,
            I => \N__5880\
        );

    \I__1181\ : CascadeMux
    port map (
            O => \N__5883\,
            I => \N__5874\
        );

    \I__1180\ : InMux
    port map (
            O => \N__5880\,
            I => \N__5871\
        );

    \I__1179\ : InMux
    port map (
            O => \N__5879\,
            I => \N__5864\
        );

    \I__1178\ : InMux
    port map (
            O => \N__5878\,
            I => \N__5864\
        );

    \I__1177\ : InMux
    port map (
            O => \N__5877\,
            I => \N__5864\
        );

    \I__1176\ : InMux
    port map (
            O => \N__5874\,
            I => \N__5861\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__5871\,
            I => \N__5856\
        );

    \I__1174\ : LocalMux
    port map (
            O => \N__5864\,
            I => \N__5856\
        );

    \I__1173\ : LocalMux
    port map (
            O => \N__5861\,
            I => \N__5853\
        );

    \I__1172\ : Span4Mux_h
    port map (
            O => \N__5856\,
            I => \N__5848\
        );

    \I__1171\ : Span4Mux_h
    port map (
            O => \N__5853\,
            I => \N__5848\
        );

    \I__1170\ : Odrv4
    port map (
            O => \N__5848\,
            I => \uut.acc_out_4\
        );

    \I__1169\ : CEMux
    port map (
            O => \N__5845\,
            I => \N__5842\
        );

    \I__1168\ : LocalMux
    port map (
            O => \N__5842\,
            I => \N__5838\
        );

    \I__1167\ : CEMux
    port map (
            O => \N__5841\,
            I => \N__5834\
        );

    \I__1166\ : Span4Mux_h
    port map (
            O => \N__5838\,
            I => \N__5830\
        );

    \I__1165\ : CEMux
    port map (
            O => \N__5837\,
            I => \N__5827\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__5834\,
            I => \N__5824\
        );

    \I__1163\ : CEMux
    port map (
            O => \N__5833\,
            I => \N__5821\
        );

    \I__1162\ : Span4Mux_v
    port map (
            O => \N__5830\,
            I => \N__5816\
        );

    \I__1161\ : LocalMux
    port map (
            O => \N__5827\,
            I => \N__5816\
        );

    \I__1160\ : Span4Mux_v
    port map (
            O => \N__5824\,
            I => \N__5813\
        );

    \I__1159\ : LocalMux
    port map (
            O => \N__5821\,
            I => \N__5810\
        );

    \I__1158\ : Span4Mux_s3_h
    port map (
            O => \N__5816\,
            I => \N__5807\
        );

    \I__1157\ : Span4Mux_h
    port map (
            O => \N__5813\,
            I => \N__5802\
        );

    \I__1156\ : Span4Mux_v
    port map (
            O => \N__5810\,
            I => \N__5802\
        );

    \I__1155\ : Odrv4
    port map (
            O => \N__5807\,
            I => \uut.ACC_LD_0_i\
        );

    \I__1154\ : Odrv4
    port map (
            O => \N__5802\,
            I => \uut.ACC_LD_0_i\
        );

    \I__1153\ : InMux
    port map (
            O => \N__5797\,
            I => \N__5794\
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__5794\,
            I => \N__5789\
        );

    \I__1151\ : InMux
    port map (
            O => \N__5793\,
            I => \N__5786\
        );

    \I__1150\ : CascadeMux
    port map (
            O => \N__5792\,
            I => \N__5783\
        );

    \I__1149\ : Span4Mux_h
    port map (
            O => \N__5789\,
            I => \N__5780\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__5786\,
            I => \N__5777\
        );

    \I__1147\ : InMux
    port map (
            O => \N__5783\,
            I => \N__5774\
        );

    \I__1146\ : Odrv4
    port map (
            O => \N__5780\,
            I => \uut.program_counter_2\
        );

    \I__1145\ : Odrv12
    port map (
            O => \N__5777\,
            I => \uut.program_counter_2\
        );

    \I__1144\ : LocalMux
    port map (
            O => \N__5774\,
            I => \uut.program_counter_2\
        );

    \I__1143\ : CascadeMux
    port map (
            O => \N__5767\,
            I => \N__5764\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5764\,
            I => \N__5760\
        );

    \I__1141\ : CascadeMux
    port map (
            O => \N__5763\,
            I => \N__5757\
        );

    \I__1140\ : LocalMux
    port map (
            O => \N__5760\,
            I => \N__5754\
        );

    \I__1139\ : InMux
    port map (
            O => \N__5757\,
            I => \N__5751\
        );

    \I__1138\ : Span4Mux_v
    port map (
            O => \N__5754\,
            I => \N__5745\
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__5751\,
            I => \N__5742\
        );

    \I__1136\ : InMux
    port map (
            O => \N__5750\,
            I => \N__5739\
        );

    \I__1135\ : CascadeMux
    port map (
            O => \N__5749\,
            I => \N__5736\
        );

    \I__1134\ : CascadeMux
    port map (
            O => \N__5748\,
            I => \N__5733\
        );

    \I__1133\ : Span4Mux_h
    port map (
            O => \N__5745\,
            I => \N__5730\
        );

    \I__1132\ : Span4Mux_s2_h
    port map (
            O => \N__5742\,
            I => \N__5725\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__5739\,
            I => \N__5725\
        );

    \I__1130\ : InMux
    port map (
            O => \N__5736\,
            I => \N__5720\
        );

    \I__1129\ : InMux
    port map (
            O => \N__5733\,
            I => \N__5720\
        );

    \I__1128\ : Odrv4
    port map (
            O => \N__5730\,
            I => \uut.program_counter_1\
        );

    \I__1127\ : Odrv4
    port map (
            O => \N__5725\,
            I => \uut.program_counter_1\
        );

    \I__1126\ : LocalMux
    port map (
            O => \N__5720\,
            I => \uut.program_counter_1\
        );

    \I__1125\ : InMux
    port map (
            O => \N__5713\,
            I => \N__5710\
        );

    \I__1124\ : LocalMux
    port map (
            O => \N__5710\,
            I => \N__5706\
        );

    \I__1123\ : InMux
    port map (
            O => \N__5709\,
            I => \N__5703\
        );

    \I__1122\ : Span4Mux_s3_h
    port map (
            O => \N__5706\,
            I => \N__5697\
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__5703\,
            I => \N__5694\
        );

    \I__1120\ : InMux
    port map (
            O => \N__5702\,
            I => \N__5687\
        );

    \I__1119\ : InMux
    port map (
            O => \N__5701\,
            I => \N__5687\
        );

    \I__1118\ : InMux
    port map (
            O => \N__5700\,
            I => \N__5687\
        );

    \I__1117\ : Odrv4
    port map (
            O => \N__5697\,
            I => \uut.program_counter_0\
        );

    \I__1116\ : Odrv12
    port map (
            O => \N__5694\,
            I => \uut.program_counter_0\
        );

    \I__1115\ : LocalMux
    port map (
            O => \N__5687\,
            I => \uut.program_counter_0\
        );

    \I__1114\ : InMux
    port map (
            O => \N__5680\,
            I => \N__5677\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__5677\,
            I => \uut.pc.program_counter_RNO_1Z0Z_2\
        );

    \I__1112\ : CascadeMux
    port map (
            O => \N__5674\,
            I => \uut.N_44_0_cascade_\
        );

    \I__1111\ : InMux
    port map (
            O => \N__5671\,
            I => \N__5668\
        );

    \I__1110\ : LocalMux
    port map (
            O => \N__5668\,
            I => \N__5665\
        );

    \I__1109\ : Odrv4
    port map (
            O => \N__5665\,
            I => \uut.pc.g0_rn_1\
        );

    \I__1108\ : CascadeMux
    port map (
            O => \N__5662\,
            I => \uut.pc.alu_out_m_0_3_cascade_\
        );

    \I__1107\ : ClkMux
    port map (
            O => \N__5659\,
            I => \N__5548\
        );

    \I__1106\ : ClkMux
    port map (
            O => \N__5658\,
            I => \N__5548\
        );

    \I__1105\ : ClkMux
    port map (
            O => \N__5657\,
            I => \N__5548\
        );

    \I__1104\ : ClkMux
    port map (
            O => \N__5656\,
            I => \N__5548\
        );

    \I__1103\ : ClkMux
    port map (
            O => \N__5655\,
            I => \N__5548\
        );

    \I__1102\ : ClkMux
    port map (
            O => \N__5654\,
            I => \N__5548\
        );

    \I__1101\ : ClkMux
    port map (
            O => \N__5653\,
            I => \N__5548\
        );

    \I__1100\ : ClkMux
    port map (
            O => \N__5652\,
            I => \N__5548\
        );

    \I__1099\ : ClkMux
    port map (
            O => \N__5651\,
            I => \N__5548\
        );

    \I__1098\ : ClkMux
    port map (
            O => \N__5650\,
            I => \N__5548\
        );

    \I__1097\ : ClkMux
    port map (
            O => \N__5649\,
            I => \N__5548\
        );

    \I__1096\ : ClkMux
    port map (
            O => \N__5648\,
            I => \N__5548\
        );

    \I__1095\ : ClkMux
    port map (
            O => \N__5647\,
            I => \N__5548\
        );

    \I__1094\ : ClkMux
    port map (
            O => \N__5646\,
            I => \N__5548\
        );

    \I__1093\ : ClkMux
    port map (
            O => \N__5645\,
            I => \N__5548\
        );

    \I__1092\ : ClkMux
    port map (
            O => \N__5644\,
            I => \N__5548\
        );

    \I__1091\ : ClkMux
    port map (
            O => \N__5643\,
            I => \N__5548\
        );

    \I__1090\ : ClkMux
    port map (
            O => \N__5642\,
            I => \N__5548\
        );

    \I__1089\ : ClkMux
    port map (
            O => \N__5641\,
            I => \N__5548\
        );

    \I__1088\ : ClkMux
    port map (
            O => \N__5640\,
            I => \N__5548\
        );

    \I__1087\ : ClkMux
    port map (
            O => \N__5639\,
            I => \N__5548\
        );

    \I__1086\ : ClkMux
    port map (
            O => \N__5638\,
            I => \N__5548\
        );

    \I__1085\ : ClkMux
    port map (
            O => \N__5637\,
            I => \N__5548\
        );

    \I__1084\ : ClkMux
    port map (
            O => \N__5636\,
            I => \N__5548\
        );

    \I__1083\ : ClkMux
    port map (
            O => \N__5635\,
            I => \N__5548\
        );

    \I__1082\ : ClkMux
    port map (
            O => \N__5634\,
            I => \N__5548\
        );

    \I__1081\ : ClkMux
    port map (
            O => \N__5633\,
            I => \N__5548\
        );

    \I__1080\ : ClkMux
    port map (
            O => \N__5632\,
            I => \N__5548\
        );

    \I__1079\ : ClkMux
    port map (
            O => \N__5631\,
            I => \N__5548\
        );

    \I__1078\ : ClkMux
    port map (
            O => \N__5630\,
            I => \N__5548\
        );

    \I__1077\ : ClkMux
    port map (
            O => \N__5629\,
            I => \N__5548\
        );

    \I__1076\ : ClkMux
    port map (
            O => \N__5628\,
            I => \N__5548\
        );

    \I__1075\ : ClkMux
    port map (
            O => \N__5627\,
            I => \N__5548\
        );

    \I__1074\ : ClkMux
    port map (
            O => \N__5626\,
            I => \N__5548\
        );

    \I__1073\ : ClkMux
    port map (
            O => \N__5625\,
            I => \N__5548\
        );

    \I__1072\ : ClkMux
    port map (
            O => \N__5624\,
            I => \N__5548\
        );

    \I__1071\ : ClkMux
    port map (
            O => \N__5623\,
            I => \N__5548\
        );

    \I__1070\ : GlobalMux
    port map (
            O => \N__5548\,
            I => \N__5545\
        );

    \I__1069\ : gio2CtrlBuf
    port map (
            O => \N__5545\,
            I => \uut.buf_clk_1_g\
        );

    \I__1068\ : CascadeMux
    port map (
            O => \N__5542\,
            I => \N__5539\
        );

    \I__1067\ : InMux
    port map (
            O => \N__5539\,
            I => \N__5536\
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__5536\,
            I => \N__5533\
        );

    \I__1065\ : Odrv4
    port map (
            O => \N__5533\,
            I => \uut.ALU_main.N_44_1\
        );

    \I__1064\ : InMux
    port map (
            O => \N__5530\,
            I => \N__5527\
        );

    \I__1063\ : LocalMux
    port map (
            O => \N__5527\,
            I => \uut.pc.g1\
        );

    \I__1062\ : CascadeMux
    port map (
            O => \N__5524\,
            I => \uut.pc.un1_inc_0_0_cascade_\
        );

    \I__1061\ : InMux
    port map (
            O => \N__5521\,
            I => \N__5517\
        );

    \I__1060\ : InMux
    port map (
            O => \N__5520\,
            I => \N__5513\
        );

    \I__1059\ : LocalMux
    port map (
            O => \N__5517\,
            I => \N__5510\
        );

    \I__1058\ : InMux
    port map (
            O => \N__5516\,
            I => \N__5507\
        );

    \I__1057\ : LocalMux
    port map (
            O => \N__5513\,
            I => \N__5502\
        );

    \I__1056\ : Span4Mux_s3_h
    port map (
            O => \N__5510\,
            I => \N__5502\
        );

    \I__1055\ : LocalMux
    port map (
            O => \N__5507\,
            I => \N__5499\
        );

    \I__1054\ : Odrv4
    port map (
            O => \N__5502\,
            I => \uut.un17_IR_OE\
        );

    \I__1053\ : Odrv12
    port map (
            O => \N__5499\,
            I => \uut.un17_IR_OE\
        );

    \I__1052\ : InMux
    port map (
            O => \N__5494\,
            I => \N__5491\
        );

    \I__1051\ : LocalMux
    port map (
            O => \N__5491\,
            I => \uut.PC_LD_0_0\
        );

    \I__1050\ : CascadeMux
    port map (
            O => \N__5488\,
            I => \uut.PC_LD_0_0_cascade_\
        );

    \I__1049\ : InMux
    port map (
            O => \N__5485\,
            I => \N__5481\
        );

    \I__1048\ : CascadeMux
    port map (
            O => \N__5484\,
            I => \N__5478\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__5481\,
            I => \N__5475\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5478\,
            I => \N__5472\
        );

    \I__1045\ : Span4Mux_v
    port map (
            O => \N__5475\,
            I => \N__5467\
        );

    \I__1044\ : LocalMux
    port map (
            O => \N__5472\,
            I => \N__5467\
        );

    \I__1043\ : Odrv4
    port map (
            O => \N__5467\,
            I => \uut.pc.un1_inc_0\
        );

    \I__1042\ : CascadeMux
    port map (
            O => \N__5464\,
            I => \uut.pc.un1_inc_0_cascade_\
        );

    \I__1041\ : InMux
    port map (
            O => \N__5461\,
            I => \N__5458\
        );

    \I__1040\ : LocalMux
    port map (
            O => \N__5458\,
            I => \N__5455\
        );

    \I__1039\ : Odrv12
    port map (
            O => \N__5455\,
            I => \uut.pc.program_counter_4_1_2\
        );

    \I__1038\ : CascadeMux
    port map (
            O => \N__5452\,
            I => \N__5448\
        );

    \I__1037\ : CascadeMux
    port map (
            O => \N__5451\,
            I => \N__5445\
        );

    \I__1036\ : InMux
    port map (
            O => \N__5448\,
            I => \N__5442\
        );

    \I__1035\ : InMux
    port map (
            O => \N__5445\,
            I => \N__5439\
        );

    \I__1034\ : LocalMux
    port map (
            O => \N__5442\,
            I => \N__5436\
        );

    \I__1033\ : LocalMux
    port map (
            O => \N__5439\,
            I => \N__5433\
        );

    \I__1032\ : Span12Mux_s10_v
    port map (
            O => \N__5436\,
            I => \N__5430\
        );

    \I__1031\ : Span4Mux_h
    port map (
            O => \N__5433\,
            I => \N__5427\
        );

    \I__1030\ : Odrv12
    port map (
            O => \N__5430\,
            I => \uut.m13\
        );

    \I__1029\ : Odrv4
    port map (
            O => \N__5427\,
            I => \uut.m13\
        );

    \I__1028\ : InMux
    port map (
            O => \N__5422\,
            I => \N__5410\
        );

    \I__1027\ : InMux
    port map (
            O => \N__5421\,
            I => \N__5407\
        );

    \I__1026\ : InMux
    port map (
            O => \N__5420\,
            I => \N__5402\
        );

    \I__1025\ : InMux
    port map (
            O => \N__5419\,
            I => \N__5402\
        );

    \I__1024\ : InMux
    port map (
            O => \N__5418\,
            I => \N__5395\
        );

    \I__1023\ : InMux
    port map (
            O => \N__5417\,
            I => \N__5395\
        );

    \I__1022\ : InMux
    port map (
            O => \N__5416\,
            I => \N__5395\
        );

    \I__1021\ : InMux
    port map (
            O => \N__5415\,
            I => \N__5388\
        );

    \I__1020\ : InMux
    port map (
            O => \N__5414\,
            I => \N__5388\
        );

    \I__1019\ : InMux
    port map (
            O => \N__5413\,
            I => \N__5388\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__5410\,
            I => \uut.q_0_fast_0\
        );

    \I__1017\ : LocalMux
    port map (
            O => \N__5407\,
            I => \uut.q_0_fast_0\
        );

    \I__1016\ : LocalMux
    port map (
            O => \N__5402\,
            I => \uut.q_0_fast_0\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__5395\,
            I => \uut.q_0_fast_0\
        );

    \I__1014\ : LocalMux
    port map (
            O => \N__5388\,
            I => \uut.q_0_fast_0\
        );

    \I__1013\ : CascadeMux
    port map (
            O => \N__5377\,
            I => \N__5373\
        );

    \I__1012\ : InMux
    port map (
            O => \N__5376\,
            I => \N__5370\
        );

    \I__1011\ : InMux
    port map (
            O => \N__5373\,
            I => \N__5367\
        );

    \I__1010\ : LocalMux
    port map (
            O => \N__5370\,
            I => \uut.seq.counter.T_fastZ0Z_2\
        );

    \I__1009\ : LocalMux
    port map (
            O => \N__5367\,
            I => \uut.seq.counter.T_fastZ0Z_2\
        );

    \I__1008\ : CascadeMux
    port map (
            O => \N__5362\,
            I => \uut.seq.counter.T_fast_RNIH09PZ0Z_2_cascade_\
        );

    \I__1007\ : InMux
    port map (
            O => \N__5359\,
            I => \N__5353\
        );

    \I__1006\ : CascadeMux
    port map (
            O => \N__5358\,
            I => \N__5350\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5357\,
            I => \N__5346\
        );

    \I__1004\ : CascadeMux
    port map (
            O => \N__5356\,
            I => \N__5343\
        );

    \I__1003\ : LocalMux
    port map (
            O => \N__5353\,
            I => \N__5336\
        );

    \I__1002\ : InMux
    port map (
            O => \N__5350\,
            I => \N__5331\
        );

    \I__1001\ : InMux
    port map (
            O => \N__5349\,
            I => \N__5331\
        );

    \I__1000\ : LocalMux
    port map (
            O => \N__5346\,
            I => \N__5328\
        );

    \I__999\ : InMux
    port map (
            O => \N__5343\,
            I => \N__5325\
        );

    \I__998\ : InMux
    port map (
            O => \N__5342\,
            I => \N__5322\
        );

    \I__997\ : InMux
    port map (
            O => \N__5341\,
            I => \N__5315\
        );

    \I__996\ : InMux
    port map (
            O => \N__5340\,
            I => \N__5315\
        );

    \I__995\ : InMux
    port map (
            O => \N__5339\,
            I => \N__5315\
        );

    \I__994\ : Odrv4
    port map (
            O => \N__5336\,
            I => \uut.ir_out_4_rep1\
        );

    \I__993\ : LocalMux
    port map (
            O => \N__5331\,
            I => \uut.ir_out_4_rep1\
        );

    \I__992\ : Odrv12
    port map (
            O => \N__5328\,
            I => \uut.ir_out_4_rep1\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__5325\,
            I => \uut.ir_out_4_rep1\
        );

    \I__990\ : LocalMux
    port map (
            O => \N__5322\,
            I => \uut.ir_out_4_rep1\
        );

    \I__989\ : LocalMux
    port map (
            O => \N__5315\,
            I => \uut.ir_out_4_rep1\
        );

    \I__988\ : InMux
    port map (
            O => \N__5302\,
            I => \N__5294\
        );

    \I__987\ : InMux
    port map (
            O => \N__5301\,
            I => \N__5289\
        );

    \I__986\ : InMux
    port map (
            O => \N__5300\,
            I => \N__5289\
        );

    \I__985\ : InMux
    port map (
            O => \N__5299\,
            I => \N__5284\
        );

    \I__984\ : InMux
    port map (
            O => \N__5298\,
            I => \N__5284\
        );

    \I__983\ : InMux
    port map (
            O => \N__5297\,
            I => \N__5280\
        );

    \I__982\ : LocalMux
    port map (
            O => \N__5294\,
            I => \N__5277\
        );

    \I__981\ : LocalMux
    port map (
            O => \N__5289\,
            I => \N__5272\
        );

    \I__980\ : LocalMux
    port map (
            O => \N__5284\,
            I => \N__5272\
        );

    \I__979\ : InMux
    port map (
            O => \N__5283\,
            I => \N__5269\
        );

    \I__978\ : LocalMux
    port map (
            O => \N__5280\,
            I => \N__5266\
        );

    \I__977\ : Span4Mux_h
    port map (
            O => \N__5277\,
            I => \N__5261\
        );

    \I__976\ : Span4Mux_v
    port map (
            O => \N__5272\,
            I => \N__5261\
        );

    \I__975\ : LocalMux
    port map (
            O => \N__5269\,
            I => \N__5258\
        );

    \I__974\ : Span4Mux_v
    port map (
            O => \N__5266\,
            I => \N__5255\
        );

    \I__973\ : Span4Mux_v
    port map (
            O => \N__5261\,
            I => \N__5250\
        );

    \I__972\ : Span4Mux_s1_v
    port map (
            O => \N__5258\,
            I => \N__5250\
        );

    \I__971\ : Odrv4
    port map (
            O => \N__5255\,
            I => \uut.ir_out_0\
        );

    \I__970\ : Odrv4
    port map (
            O => \N__5250\,
            I => \uut.ir_out_0\
        );

    \I__969\ : CascadeMux
    port map (
            O => \N__5245\,
            I => \N__5238\
        );

    \I__968\ : InMux
    port map (
            O => \N__5244\,
            I => \N__5234\
        );

    \I__967\ : InMux
    port map (
            O => \N__5243\,
            I => \N__5231\
        );

    \I__966\ : InMux
    port map (
            O => \N__5242\,
            I => \N__5226\
        );

    \I__965\ : InMux
    port map (
            O => \N__5241\,
            I => \N__5226\
        );

    \I__964\ : InMux
    port map (
            O => \N__5238\,
            I => \N__5221\
        );

    \I__963\ : InMux
    port map (
            O => \N__5237\,
            I => \N__5221\
        );

    \I__962\ : LocalMux
    port map (
            O => \N__5234\,
            I => \N__5214\
        );

    \I__961\ : LocalMux
    port map (
            O => \N__5231\,
            I => \N__5214\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__5226\,
            I => \N__5214\
        );

    \I__959\ : LocalMux
    port map (
            O => \N__5221\,
            I => \uut.acc_out_0\
        );

    \I__958\ : Odrv12
    port map (
            O => \N__5214\,
            I => \uut.acc_out_0\
        );

    \I__957\ : CascadeMux
    port map (
            O => \N__5209\,
            I => \uut.OUT_LD_cascade_\
        );

    \I__956\ : InMux
    port map (
            O => \N__5206\,
            I => \N__5203\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__5203\,
            I => \N__5200\
        );

    \I__954\ : Span4Mux_v
    port map (
            O => \N__5200\,
            I => \N__5197\
        );

    \I__953\ : Odrv4
    port map (
            O => \N__5197\,
            I => \uut.pc.G_26_i_a4_1\
        );

    \I__952\ : CascadeMux
    port map (
            O => \N__5194\,
            I => \N__5189\
        );

    \I__951\ : CascadeMux
    port map (
            O => \N__5193\,
            I => \N__5186\
        );

    \I__950\ : CascadeMux
    port map (
            O => \N__5192\,
            I => \N__5183\
        );

    \I__949\ : InMux
    port map (
            O => \N__5189\,
            I => \N__5178\
        );

    \I__948\ : InMux
    port map (
            O => \N__5186\,
            I => \N__5175\
        );

    \I__947\ : InMux
    port map (
            O => \N__5183\,
            I => \N__5172\
        );

    \I__946\ : InMux
    port map (
            O => \N__5182\,
            I => \N__5168\
        );

    \I__945\ : InMux
    port map (
            O => \N__5181\,
            I => \N__5165\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__5178\,
            I => \N__5160\
        );

    \I__943\ : LocalMux
    port map (
            O => \N__5175\,
            I => \N__5160\
        );

    \I__942\ : LocalMux
    port map (
            O => \N__5172\,
            I => \N__5157\
        );

    \I__941\ : InMux
    port map (
            O => \N__5171\,
            I => \N__5154\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__5168\,
            I => \N__5149\
        );

    \I__939\ : LocalMux
    port map (
            O => \N__5165\,
            I => \N__5149\
        );

    \I__938\ : Span4Mux_v
    port map (
            O => \N__5160\,
            I => \N__5146\
        );

    \I__937\ : Span4Mux_h
    port map (
            O => \N__5157\,
            I => \N__5143\
        );

    \I__936\ : LocalMux
    port map (
            O => \N__5154\,
            I => \uut.acc_out_1\
        );

    \I__935\ : Odrv12
    port map (
            O => \N__5149\,
            I => \uut.acc_out_1\
        );

    \I__934\ : Odrv4
    port map (
            O => \N__5146\,
            I => \uut.acc_out_1\
        );

    \I__933\ : Odrv4
    port map (
            O => \N__5143\,
            I => \uut.acc_out_1\
        );

    \I__932\ : CascadeMux
    port map (
            O => \N__5134\,
            I => \uut.ALU_main.ALU_Out_0Z0Z_1_cascade_\
        );

    \I__931\ : InMux
    port map (
            O => \N__5131\,
            I => \N__5128\
        );

    \I__930\ : LocalMux
    port map (
            O => \N__5128\,
            I => \N__5125\
        );

    \I__929\ : Span4Mux_s2_h
    port map (
            O => \N__5125\,
            I => \N__5121\
        );

    \I__928\ : InMux
    port map (
            O => \N__5124\,
            I => \N__5118\
        );

    \I__927\ : Odrv4
    port map (
            O => \N__5121\,
            I => \uut.un1_A_cry_0_c_RNI3CH45\
        );

    \I__926\ : LocalMux
    port map (
            O => \N__5118\,
            I => \uut.un1_A_cry_0_c_RNI3CH45\
        );

    \I__925\ : InMux
    port map (
            O => \N__5113\,
            I => \N__5110\
        );

    \I__924\ : LocalMux
    port map (
            O => \N__5110\,
            I => \N__5107\
        );

    \I__923\ : Span4Mux_v
    port map (
            O => \N__5107\,
            I => \N__5104\
        );

    \I__922\ : Odrv4
    port map (
            O => \N__5104\,
            I => \uut.seq.counter.un2_MAR_LD\
        );

    \I__921\ : InMux
    port map (
            O => \N__5101\,
            I => \N__5096\
        );

    \I__920\ : CascadeMux
    port map (
            O => \N__5100\,
            I => \N__5093\
        );

    \I__919\ : InMux
    port map (
            O => \N__5099\,
            I => \N__5089\
        );

    \I__918\ : LocalMux
    port map (
            O => \N__5096\,
            I => \N__5086\
        );

    \I__917\ : InMux
    port map (
            O => \N__5093\,
            I => \N__5083\
        );

    \I__916\ : CascadeMux
    port map (
            O => \N__5092\,
            I => \N__5077\
        );

    \I__915\ : LocalMux
    port map (
            O => \N__5089\,
            I => \N__5074\
        );

    \I__914\ : Span4Mux_v
    port map (
            O => \N__5086\,
            I => \N__5069\
        );

    \I__913\ : LocalMux
    port map (
            O => \N__5083\,
            I => \N__5069\
        );

    \I__912\ : InMux
    port map (
            O => \N__5082\,
            I => \N__5064\
        );

    \I__911\ : InMux
    port map (
            O => \N__5081\,
            I => \N__5064\
        );

    \I__910\ : InMux
    port map (
            O => \N__5080\,
            I => \N__5061\
        );

    \I__909\ : InMux
    port map (
            O => \N__5077\,
            I => \N__5058\
        );

    \I__908\ : Odrv12
    port map (
            O => \N__5074\,
            I => \uut.T_2_rep1\
        );

    \I__907\ : Odrv4
    port map (
            O => \N__5069\,
            I => \uut.T_2_rep1\
        );

    \I__906\ : LocalMux
    port map (
            O => \N__5064\,
            I => \uut.T_2_rep1\
        );

    \I__905\ : LocalMux
    port map (
            O => \N__5061\,
            I => \uut.T_2_rep1\
        );

    \I__904\ : LocalMux
    port map (
            O => \N__5058\,
            I => \uut.T_2_rep1\
        );

    \I__903\ : InMux
    port map (
            O => \N__5047\,
            I => \N__5044\
        );

    \I__902\ : LocalMux
    port map (
            O => \N__5044\,
            I => \uut.seq.counter.T_2_rep1_RNIV9NUZ0\
        );

    \I__901\ : InMux
    port map (
            O => \N__5041\,
            I => \N__5038\
        );

    \I__900\ : LocalMux
    port map (
            O => \N__5038\,
            I => \N__5035\
        );

    \I__899\ : Span4Mux_h
    port map (
            O => \N__5035\,
            I => \N__5032\
        );

    \I__898\ : Odrv4
    port map (
            O => \N__5032\,
            I => \uut.bus_5\
        );

    \I__897\ : CascadeMux
    port map (
            O => \N__5029\,
            I => \N__5025\
        );

    \I__896\ : CascadeMux
    port map (
            O => \N__5028\,
            I => \N__5022\
        );

    \I__895\ : InMux
    port map (
            O => \N__5025\,
            I => \N__5016\
        );

    \I__894\ : InMux
    port map (
            O => \N__5022\,
            I => \N__5016\
        );

    \I__893\ : CascadeMux
    port map (
            O => \N__5021\,
            I => \N__5013\
        );

    \I__892\ : LocalMux
    port map (
            O => \N__5016\,
            I => \N__5009\
        );

    \I__891\ : InMux
    port map (
            O => \N__5013\,
            I => \N__5006\
        );

    \I__890\ : InMux
    port map (
            O => \N__5012\,
            I => \N__5003\
        );

    \I__889\ : Odrv4
    port map (
            O => \N__5009\,
            I => \uut.q_0_fast_1\
        );

    \I__888\ : LocalMux
    port map (
            O => \N__5006\,
            I => \uut.q_0_fast_1\
        );

    \I__887\ : LocalMux
    port map (
            O => \N__5003\,
            I => \uut.q_0_fast_1\
        );

    \I__886\ : InMux
    port map (
            O => \N__4996\,
            I => \N__4993\
        );

    \I__885\ : LocalMux
    port map (
            O => \N__4993\,
            I => \uut.seq.counter.T_1_fastZ0Z_0\
        );

    \I__884\ : InMux
    port map (
            O => \N__4990\,
            I => \N__4983\
        );

    \I__883\ : InMux
    port map (
            O => \N__4989\,
            I => \N__4983\
        );

    \I__882\ : CascadeMux
    port map (
            O => \N__4988\,
            I => \N__4974\
        );

    \I__881\ : LocalMux
    port map (
            O => \N__4983\,
            I => \N__4971\
        );

    \I__880\ : InMux
    port map (
            O => \N__4982\,
            I => \N__4968\
        );

    \I__879\ : InMux
    port map (
            O => \N__4981\,
            I => \N__4965\
        );

    \I__878\ : InMux
    port map (
            O => \N__4980\,
            I => \N__4962\
        );

    \I__877\ : InMux
    port map (
            O => \N__4979\,
            I => \N__4959\
        );

    \I__876\ : InMux
    port map (
            O => \N__4978\,
            I => \N__4954\
        );

    \I__875\ : InMux
    port map (
            O => \N__4977\,
            I => \N__4954\
        );

    \I__874\ : InMux
    port map (
            O => \N__4974\,
            I => \N__4951\
        );

    \I__873\ : Odrv12
    port map (
            O => \N__4971\,
            I => \uut.ir_out_fast_4\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__4968\,
            I => \uut.ir_out_fast_4\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__4965\,
            I => \uut.ir_out_fast_4\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__4962\,
            I => \uut.ir_out_fast_4\
        );

    \I__869\ : LocalMux
    port map (
            O => \N__4959\,
            I => \uut.ir_out_fast_4\
        );

    \I__868\ : LocalMux
    port map (
            O => \N__4954\,
            I => \uut.ir_out_fast_4\
        );

    \I__867\ : LocalMux
    port map (
            O => \N__4951\,
            I => \uut.ir_out_fast_4\
        );

    \I__866\ : InMux
    port map (
            O => \N__4936\,
            I => \N__4933\
        );

    \I__865\ : LocalMux
    port map (
            O => \N__4933\,
            I => \N__4925\
        );

    \I__864\ : InMux
    port map (
            O => \N__4932\,
            I => \N__4922\
        );

    \I__863\ : InMux
    port map (
            O => \N__4931\,
            I => \N__4917\
        );

    \I__862\ : InMux
    port map (
            O => \N__4930\,
            I => \N__4917\
        );

    \I__861\ : InMux
    port map (
            O => \N__4929\,
            I => \N__4914\
        );

    \I__860\ : InMux
    port map (
            O => \N__4928\,
            I => \N__4911\
        );

    \I__859\ : Span4Mux_h
    port map (
            O => \N__4925\,
            I => \N__4901\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__4922\,
            I => \N__4901\
        );

    \I__857\ : LocalMux
    port map (
            O => \N__4917\,
            I => \N__4898\
        );

    \I__856\ : LocalMux
    port map (
            O => \N__4914\,
            I => \N__4893\
        );

    \I__855\ : LocalMux
    port map (
            O => \N__4911\,
            I => \N__4893\
        );

    \I__854\ : InMux
    port map (
            O => \N__4910\,
            I => \N__4888\
        );

    \I__853\ : InMux
    port map (
            O => \N__4909\,
            I => \N__4888\
        );

    \I__852\ : InMux
    port map (
            O => \N__4908\,
            I => \N__4881\
        );

    \I__851\ : InMux
    port map (
            O => \N__4907\,
            I => \N__4881\
        );

    \I__850\ : InMux
    port map (
            O => \N__4906\,
            I => \N__4881\
        );

    \I__849\ : Odrv4
    port map (
            O => \N__4901\,
            I => \uut.ir_out_5\
        );

    \I__848\ : Odrv12
    port map (
            O => \N__4898\,
            I => \uut.ir_out_5\
        );

    \I__847\ : Odrv4
    port map (
            O => \N__4893\,
            I => \uut.ir_out_5\
        );

    \I__846\ : LocalMux
    port map (
            O => \N__4888\,
            I => \uut.ir_out_5\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__4881\,
            I => \uut.ir_out_5\
        );

    \I__844\ : InMux
    port map (
            O => \N__4870\,
            I => \N__4866\
        );

    \I__843\ : InMux
    port map (
            O => \N__4869\,
            I => \N__4860\
        );

    \I__842\ : LocalMux
    port map (
            O => \N__4866\,
            I => \N__4857\
        );

    \I__841\ : InMux
    port map (
            O => \N__4865\,
            I => \N__4850\
        );

    \I__840\ : InMux
    port map (
            O => \N__4864\,
            I => \N__4850\
        );

    \I__839\ : InMux
    port map (
            O => \N__4863\,
            I => \N__4850\
        );

    \I__838\ : LocalMux
    port map (
            O => \N__4860\,
            I => \uut.q_ret_1_fast\
        );

    \I__837\ : Odrv4
    port map (
            O => \N__4857\,
            I => \uut.q_ret_1_fast\
        );

    \I__836\ : LocalMux
    port map (
            O => \N__4850\,
            I => \uut.q_ret_1_fast\
        );

    \I__835\ : InMux
    port map (
            O => \N__4843\,
            I => \N__4836\
        );

    \I__834\ : InMux
    port map (
            O => \N__4842\,
            I => \N__4833\
        );

    \I__833\ : InMux
    port map (
            O => \N__4841\,
            I => \N__4830\
        );

    \I__832\ : InMux
    port map (
            O => \N__4840\,
            I => \N__4827\
        );

    \I__831\ : InMux
    port map (
            O => \N__4839\,
            I => \N__4824\
        );

    \I__830\ : LocalMux
    port map (
            O => \N__4836\,
            I => \uut.seq.counter.T_4\
        );

    \I__829\ : LocalMux
    port map (
            O => \N__4833\,
            I => \uut.seq.counter.T_4\
        );

    \I__828\ : LocalMux
    port map (
            O => \N__4830\,
            I => \uut.seq.counter.T_4\
        );

    \I__827\ : LocalMux
    port map (
            O => \N__4827\,
            I => \uut.seq.counter.T_4\
        );

    \I__826\ : LocalMux
    port map (
            O => \N__4824\,
            I => \uut.seq.counter.T_4\
        );

    \I__825\ : CascadeMux
    port map (
            O => \N__4813\,
            I => \uut.seq.un10_ACC_LD_xZ0Z1_cascade_\
        );

    \I__824\ : CascadeMux
    port map (
            O => \N__4810\,
            I => \uut.T_1_fast_RNI28LI1_0_cascade_\
        );

    \I__823\ : InMux
    port map (
            O => \N__4807\,
            I => \N__4800\
        );

    \I__822\ : InMux
    port map (
            O => \N__4806\,
            I => \N__4800\
        );

    \I__821\ : InMux
    port map (
            O => \N__4805\,
            I => \N__4797\
        );

    \I__820\ : LocalMux
    port map (
            O => \N__4800\,
            I => \N__4792\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__4797\,
            I => \N__4792\
        );

    \I__818\ : Span4Mux_v
    port map (
            O => \N__4792\,
            I => \N__4789\
        );

    \I__817\ : Odrv4
    port map (
            O => \N__4789\,
            I => \uut.N_41\
        );

    \I__816\ : CascadeMux
    port map (
            O => \N__4786\,
            I => \uut.seq.counter.T_2_rep1_RNIJDGJZ0_cascade_\
        );

    \I__815\ : InMux
    port map (
            O => \N__4783\,
            I => \N__4779\
        );

    \I__814\ : InMux
    port map (
            O => \N__4782\,
            I => \N__4776\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__4779\,
            I => \uut.seq.D_4\
        );

    \I__812\ : LocalMux
    port map (
            O => \N__4776\,
            I => \uut.seq.D_4\
        );

    \I__811\ : CascadeMux
    port map (
            O => \N__4771\,
            I => \uut.D_1_3_cascade_\
        );

    \I__810\ : InMux
    port map (
            O => \N__4768\,
            I => \N__4764\
        );

    \I__809\ : InMux
    port map (
            O => \N__4767\,
            I => \N__4761\
        );

    \I__808\ : LocalMux
    port map (
            O => \N__4764\,
            I => \N__4754\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__4761\,
            I => \N__4751\
        );

    \I__806\ : InMux
    port map (
            O => \N__4760\,
            I => \N__4746\
        );

    \I__805\ : InMux
    port map (
            O => \N__4759\,
            I => \N__4746\
        );

    \I__804\ : CascadeMux
    port map (
            O => \N__4758\,
            I => \N__4743\
        );

    \I__803\ : CascadeMux
    port map (
            O => \N__4757\,
            I => \N__4740\
        );

    \I__802\ : Span4Mux_h
    port map (
            O => \N__4754\,
            I => \N__4733\
        );

    \I__801\ : Span4Mux_h
    port map (
            O => \N__4751\,
            I => \N__4730\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__4746\,
            I => \N__4727\
        );

    \I__799\ : InMux
    port map (
            O => \N__4743\,
            I => \N__4714\
        );

    \I__798\ : InMux
    port map (
            O => \N__4740\,
            I => \N__4714\
        );

    \I__797\ : InMux
    port map (
            O => \N__4739\,
            I => \N__4714\
        );

    \I__796\ : InMux
    port map (
            O => \N__4738\,
            I => \N__4714\
        );

    \I__795\ : InMux
    port map (
            O => \N__4737\,
            I => \N__4714\
        );

    \I__794\ : InMux
    port map (
            O => \N__4736\,
            I => \N__4714\
        );

    \I__793\ : Odrv4
    port map (
            O => \N__4733\,
            I => \uut.un7_ACC_LD\
        );

    \I__792\ : Odrv4
    port map (
            O => \N__4730\,
            I => \uut.un7_ACC_LD\
        );

    \I__791\ : Odrv4
    port map (
            O => \N__4727\,
            I => \uut.un7_ACC_LD\
        );

    \I__790\ : LocalMux
    port map (
            O => \N__4714\,
            I => \uut.un7_ACC_LD\
        );

    \I__789\ : InMux
    port map (
            O => \N__4705\,
            I => \N__4697\
        );

    \I__788\ : InMux
    port map (
            O => \N__4704\,
            I => \N__4692\
        );

    \I__787\ : InMux
    port map (
            O => \N__4703\,
            I => \N__4692\
        );

    \I__786\ : InMux
    port map (
            O => \N__4702\,
            I => \N__4689\
        );

    \I__785\ : InMux
    port map (
            O => \N__4701\,
            I => \N__4686\
        );

    \I__784\ : InMux
    port map (
            O => \N__4700\,
            I => \N__4681\
        );

    \I__783\ : LocalMux
    port map (
            O => \N__4697\,
            I => \N__4678\
        );

    \I__782\ : LocalMux
    port map (
            O => \N__4692\,
            I => \N__4674\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__4689\,
            I => \N__4671\
        );

    \I__780\ : LocalMux
    port map (
            O => \N__4686\,
            I => \N__4668\
        );

    \I__779\ : InMux
    port map (
            O => \N__4685\,
            I => \N__4663\
        );

    \I__778\ : InMux
    port map (
            O => \N__4684\,
            I => \N__4663\
        );

    \I__777\ : LocalMux
    port map (
            O => \N__4681\,
            I => \N__4658\
        );

    \I__776\ : Span4Mux_h
    port map (
            O => \N__4678\,
            I => \N__4658\
        );

    \I__775\ : InMux
    port map (
            O => \N__4677\,
            I => \N__4655\
        );

    \I__774\ : Odrv4
    port map (
            O => \N__4674\,
            I => \uut.ir_out_4\
        );

    \I__773\ : Odrv4
    port map (
            O => \N__4671\,
            I => \uut.ir_out_4\
        );

    \I__772\ : Odrv12
    port map (
            O => \N__4668\,
            I => \uut.ir_out_4\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__4663\,
            I => \uut.ir_out_4\
        );

    \I__770\ : Odrv4
    port map (
            O => \N__4658\,
            I => \uut.ir_out_4\
        );

    \I__769\ : LocalMux
    port map (
            O => \N__4655\,
            I => \uut.ir_out_4\
        );

    \I__768\ : InMux
    port map (
            O => \N__4642\,
            I => \N__4638\
        );

    \I__767\ : InMux
    port map (
            O => \N__4641\,
            I => \N__4635\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__4638\,
            I => \uut.seq.counter.T_1_fastZ0Z_3\
        );

    \I__765\ : LocalMux
    port map (
            O => \N__4635\,
            I => \uut.seq.counter.T_1_fastZ0Z_3\
        );

    \I__764\ : CascadeMux
    port map (
            O => \N__4630\,
            I => \uut.seq.counter.T_4_cascade_\
        );

    \I__763\ : InMux
    port map (
            O => \N__4627\,
            I => \N__4624\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__4624\,
            I => \N__4621\
        );

    \I__761\ : Span4Mux_s3_h
    port map (
            O => \N__4621\,
            I => \N__4618\
        );

    \I__760\ : Odrv4
    port map (
            O => \N__4618\,
            I => \uut.seq.counter.T_1_fast_RNI4JTR1_0Z0Z_0\
        );

    \I__759\ : InMux
    port map (
            O => \N__4615\,
            I => \N__4612\
        );

    \I__758\ : LocalMux
    port map (
            O => \N__4612\,
            I => \N__4609\
        );

    \I__757\ : Span4Mux_h
    port map (
            O => \N__4609\,
            I => \N__4606\
        );

    \I__756\ : Odrv4
    port map (
            O => \N__4606\,
            I => \uut.ALU_main.un1_A_cry_5_c_RNINKZ0Z655\
        );

    \I__755\ : InMux
    port map (
            O => \N__4603\,
            I => \uut.ALU_main.un1_A_cry_5\
        );

    \I__754\ : InMux
    port map (
            O => \N__4600\,
            I => \bfn_9_13_0_\
        );

    \I__753\ : InMux
    port map (
            O => \N__4597\,
            I => \N__4594\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__4594\,
            I => \N__4591\
        );

    \I__751\ : Odrv12
    port map (
            O => \N__4591\,
            I => \uut.ALU_main.un1_A_cry_6_c_RNINIMNZ0Z4\
        );

    \I__750\ : InMux
    port map (
            O => \N__4588\,
            I => \N__4585\
        );

    \I__749\ : LocalMux
    port map (
            O => \N__4585\,
            I => \uut.ALU_main.un1_A_axb_1_l_ofxZ0\
        );

    \I__748\ : InMux
    port map (
            O => \N__4582\,
            I => \N__4578\
        );

    \I__747\ : InMux
    port map (
            O => \N__4581\,
            I => \N__4575\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__4578\,
            I => \N__4572\
        );

    \I__745\ : LocalMux
    port map (
            O => \N__4575\,
            I => \N__4569\
        );

    \I__744\ : Odrv4
    port map (
            O => \N__4572\,
            I => \uut.b_reg_out_6\
        );

    \I__743\ : Odrv12
    port map (
            O => \N__4569\,
            I => \uut.b_reg_out_6\
        );

    \I__742\ : InMux
    port map (
            O => \N__4564\,
            I => \N__4561\
        );

    \I__741\ : LocalMux
    port map (
            O => \N__4561\,
            I => \uut.ALU_main.un1_A_axb_6_l_ofxZ0\
        );

    \I__740\ : InMux
    port map (
            O => \N__4558\,
            I => \N__4555\
        );

    \I__739\ : LocalMux
    port map (
            O => \N__4555\,
            I => \N__4551\
        );

    \I__738\ : InMux
    port map (
            O => \N__4554\,
            I => \N__4548\
        );

    \I__737\ : Span4Mux_h
    port map (
            O => \N__4551\,
            I => \N__4545\
        );

    \I__736\ : LocalMux
    port map (
            O => \N__4548\,
            I => \uut.b_reg_out_5\
        );

    \I__735\ : Odrv4
    port map (
            O => \N__4545\,
            I => \uut.b_reg_out_5\
        );

    \I__734\ : InMux
    port map (
            O => \N__4540\,
            I => \N__4537\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__4537\,
            I => \uut.ALU_main.un1_A_axb_5_l_ofxZ0\
        );

    \I__732\ : CascadeMux
    port map (
            O => \N__4534\,
            I => \N__4531\
        );

    \I__731\ : InMux
    port map (
            O => \N__4531\,
            I => \N__4528\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__4528\,
            I => \uut.ALU_main.un1_A_axb_0_l_ofxZ0\
        );

    \I__729\ : InMux
    port map (
            O => \N__4525\,
            I => \N__4521\
        );

    \I__728\ : InMux
    port map (
            O => \N__4524\,
            I => \N__4518\
        );

    \I__727\ : LocalMux
    port map (
            O => \N__4521\,
            I => \N__4515\
        );

    \I__726\ : LocalMux
    port map (
            O => \N__4518\,
            I => \uut.b_reg_out_7\
        );

    \I__725\ : Odrv12
    port map (
            O => \N__4515\,
            I => \uut.b_reg_out_7\
        );

    \I__724\ : InMux
    port map (
            O => \N__4510\,
            I => \N__4507\
        );

    \I__723\ : LocalMux
    port map (
            O => \N__4507\,
            I => \uut.ALU_main.un1_A_axbZ0Z_7\
        );

    \I__722\ : InMux
    port map (
            O => \N__4504\,
            I => \N__4501\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__4501\,
            I => \N__4496\
        );

    \I__720\ : InMux
    port map (
            O => \N__4500\,
            I => \N__4493\
        );

    \I__719\ : InMux
    port map (
            O => \N__4499\,
            I => \N__4490\
        );

    \I__718\ : Span4Mux_h
    port map (
            O => \N__4496\,
            I => \N__4487\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__4493\,
            I => \uut.b_reg_out_2\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__4490\,
            I => \uut.b_reg_out_2\
        );

    \I__715\ : Odrv4
    port map (
            O => \N__4487\,
            I => \uut.b_reg_out_2\
        );

    \I__714\ : CascadeMux
    port map (
            O => \N__4480\,
            I => \N__4475\
        );

    \I__713\ : CascadeMux
    port map (
            O => \N__4479\,
            I => \N__4472\
        );

    \I__712\ : InMux
    port map (
            O => \N__4478\,
            I => \N__4469\
        );

    \I__711\ : InMux
    port map (
            O => \N__4475\,
            I => \N__4463\
        );

    \I__710\ : InMux
    port map (
            O => \N__4472\,
            I => \N__4460\
        );

    \I__709\ : LocalMux
    port map (
            O => \N__4469\,
            I => \N__4457\
        );

    \I__708\ : InMux
    port map (
            O => \N__4468\,
            I => \N__4454\
        );

    \I__707\ : InMux
    port map (
            O => \N__4467\,
            I => \N__4451\
        );

    \I__706\ : InMux
    port map (
            O => \N__4466\,
            I => \N__4448\
        );

    \I__705\ : LocalMux
    port map (
            O => \N__4463\,
            I => \N__4443\
        );

    \I__704\ : LocalMux
    port map (
            O => \N__4460\,
            I => \N__4443\
        );

    \I__703\ : Span4Mux_v
    port map (
            O => \N__4457\,
            I => \N__4438\
        );

    \I__702\ : LocalMux
    port map (
            O => \N__4454\,
            I => \N__4438\
        );

    \I__701\ : LocalMux
    port map (
            O => \N__4451\,
            I => \N__4435\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__4448\,
            I => \N__4430\
        );

    \I__699\ : Span4Mux_v
    port map (
            O => \N__4443\,
            I => \N__4430\
        );

    \I__698\ : Odrv4
    port map (
            O => \N__4438\,
            I => \uut.acc_out_2\
        );

    \I__697\ : Odrv4
    port map (
            O => \N__4435\,
            I => \uut.acc_out_2\
        );

    \I__696\ : Odrv4
    port map (
            O => \N__4430\,
            I => \uut.acc_out_2\
        );

    \I__695\ : InMux
    port map (
            O => \N__4423\,
            I => \N__4420\
        );

    \I__694\ : LocalMux
    port map (
            O => \N__4420\,
            I => \N__4412\
        );

    \I__693\ : InMux
    port map (
            O => \N__4419\,
            I => \N__4409\
        );

    \I__692\ : InMux
    port map (
            O => \N__4418\,
            I => \N__4406\
        );

    \I__691\ : InMux
    port map (
            O => \N__4417\,
            I => \N__4401\
        );

    \I__690\ : InMux
    port map (
            O => \N__4416\,
            I => \N__4401\
        );

    \I__689\ : CascadeMux
    port map (
            O => \N__4415\,
            I => \N__4393\
        );

    \I__688\ : Span4Mux_v
    port map (
            O => \N__4412\,
            I => \N__4390\
        );

    \I__687\ : LocalMux
    port map (
            O => \N__4409\,
            I => \N__4385\
        );

    \I__686\ : LocalMux
    port map (
            O => \N__4406\,
            I => \N__4385\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__4401\,
            I => \N__4382\
        );

    \I__684\ : InMux
    port map (
            O => \N__4400\,
            I => \N__4371\
        );

    \I__683\ : InMux
    port map (
            O => \N__4399\,
            I => \N__4371\
        );

    \I__682\ : InMux
    port map (
            O => \N__4398\,
            I => \N__4371\
        );

    \I__681\ : InMux
    port map (
            O => \N__4397\,
            I => \N__4371\
        );

    \I__680\ : InMux
    port map (
            O => \N__4396\,
            I => \N__4371\
        );

    \I__679\ : InMux
    port map (
            O => \N__4393\,
            I => \N__4368\
        );

    \I__678\ : Odrv4
    port map (
            O => \N__4390\,
            I => \uut.un13_ACC_LD\
        );

    \I__677\ : Odrv4
    port map (
            O => \N__4385\,
            I => \uut.un13_ACC_LD\
        );

    \I__676\ : Odrv4
    port map (
            O => \N__4382\,
            I => \uut.un13_ACC_LD\
        );

    \I__675\ : LocalMux
    port map (
            O => \N__4371\,
            I => \uut.un13_ACC_LD\
        );

    \I__674\ : LocalMux
    port map (
            O => \N__4368\,
            I => \uut.un13_ACC_LD\
        );

    \I__673\ : InMux
    port map (
            O => \N__4357\,
            I => \N__4354\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__4354\,
            I => \uut.ALU_main.un1_A_axb_2_l_ofxZ0\
        );

    \I__671\ : InMux
    port map (
            O => \N__4351\,
            I => \N__4348\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__4348\,
            I => \uut.pc.program_counter_0_1_1\
        );

    \I__669\ : CascadeMux
    port map (
            O => \N__4345\,
            I => \N__4342\
        );

    \I__668\ : InMux
    port map (
            O => \N__4342\,
            I => \N__4338\
        );

    \I__667\ : InMux
    port map (
            O => \N__4341\,
            I => \N__4335\
        );

    \I__666\ : LocalMux
    port map (
            O => \N__4338\,
            I => \N__4330\
        );

    \I__665\ : LocalMux
    port map (
            O => \N__4335\,
            I => \N__4330\
        );

    \I__664\ : Odrv4
    port map (
            O => \N__4330\,
            I => \uut.S0_0_i\
        );

    \I__663\ : InMux
    port map (
            O => \N__4327\,
            I => \N__4321\
        );

    \I__662\ : InMux
    port map (
            O => \N__4326\,
            I => \N__4321\
        );

    \I__661\ : LocalMux
    port map (
            O => \N__4321\,
            I => \N__4317\
        );

    \I__660\ : InMux
    port map (
            O => \N__4320\,
            I => \N__4314\
        );

    \I__659\ : Odrv4
    port map (
            O => \N__4317\,
            I => \uut.un1_A_cry_0_s\
        );

    \I__658\ : LocalMux
    port map (
            O => \N__4314\,
            I => \uut.un1_A_cry_0_s\
        );

    \I__657\ : InMux
    port map (
            O => \N__4309\,
            I => \uut.ALU_main.un1_A_cry_0_c_THRU_CO\
        );

    \I__656\ : InMux
    port map (
            O => \N__4306\,
            I => \uut.ALU_main.un1_A_cry_0\
        );

    \I__655\ : InMux
    port map (
            O => \N__4303\,
            I => \N__4300\
        );

    \I__654\ : LocalMux
    port map (
            O => \N__4300\,
            I => \N__4297\
        );

    \I__653\ : Span4Mux_v
    port map (
            O => \N__4297\,
            I => \N__4293\
        );

    \I__652\ : InMux
    port map (
            O => \N__4296\,
            I => \N__4290\
        );

    \I__651\ : Odrv4
    port map (
            O => \N__4293\,
            I => \uut.ALU_main.un1_A_cry_1_c_RNI7KLZ0Z45\
        );

    \I__650\ : LocalMux
    port map (
            O => \N__4290\,
            I => \uut.ALU_main.un1_A_cry_1_c_RNI7KLZ0Z45\
        );

    \I__649\ : InMux
    port map (
            O => \N__4285\,
            I => \uut.ALU_main.un1_A_cry_1\
        );

    \I__648\ : InMux
    port map (
            O => \N__4282\,
            I => \N__4279\
        );

    \I__647\ : LocalMux
    port map (
            O => \N__4279\,
            I => \uut.ALU_main.un1_A_axb_3_l_ofxZ0\
        );

    \I__646\ : InMux
    port map (
            O => \N__4276\,
            I => \uut.ALU_main.un1_A_cry_2_cZ0\
        );

    \I__645\ : InMux
    port map (
            O => \N__4273\,
            I => \N__4270\
        );

    \I__644\ : LocalMux
    port map (
            O => \N__4270\,
            I => \N__4267\
        );

    \I__643\ : Odrv4
    port map (
            O => \N__4267\,
            I => \uut.ALU_main.un1_A_axb_4_l_ofxZ0\
        );

    \I__642\ : InMux
    port map (
            O => \N__4264\,
            I => \N__4261\
        );

    \I__641\ : LocalMux
    port map (
            O => \N__4261\,
            I => \N__4258\
        );

    \I__640\ : Odrv4
    port map (
            O => \N__4258\,
            I => \uut.ALU_main.un1_A_cry_3_c_RNIF4UZ0Z45\
        );

    \I__639\ : InMux
    port map (
            O => \N__4255\,
            I => \uut.ALU_main.un1_A_cry_3\
        );

    \I__638\ : InMux
    port map (
            O => \N__4252\,
            I => \N__4249\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__4249\,
            I => \N__4246\
        );

    \I__636\ : Odrv4
    port map (
            O => \N__4246\,
            I => \uut.ALU_main.un1_A_cry_4_c_RNIJCZ0Z255\
        );

    \I__635\ : InMux
    port map (
            O => \N__4243\,
            I => \uut.ALU_main.un1_A_cry_4\
        );

    \I__634\ : InMux
    port map (
            O => \N__4240\,
            I => \N__4236\
        );

    \I__633\ : InMux
    port map (
            O => \N__4239\,
            I => \N__4233\
        );

    \I__632\ : LocalMux
    port map (
            O => \N__4236\,
            I => \N__4228\
        );

    \I__631\ : LocalMux
    port map (
            O => \N__4233\,
            I => \N__4228\
        );

    \I__630\ : Odrv4
    port map (
            O => \N__4228\,
            I => \uut.T_1_RNIVVKI3_3\
        );

    \I__629\ : InMux
    port map (
            O => \N__4225\,
            I => \N__4220\
        );

    \I__628\ : InMux
    port map (
            O => \N__4224\,
            I => \N__4215\
        );

    \I__627\ : InMux
    port map (
            O => \N__4223\,
            I => \N__4215\
        );

    \I__626\ : LocalMux
    port map (
            O => \N__4220\,
            I => \uut.program_counter_m_0\
        );

    \I__625\ : LocalMux
    port map (
            O => \N__4215\,
            I => \uut.program_counter_m_0\
        );

    \I__624\ : CascadeMux
    port map (
            O => \N__4210\,
            I => \uut.pc.G_26_i_a4_5_sx_cascade_\
        );

    \I__623\ : InMux
    port map (
            O => \N__4207\,
            I => \N__4204\
        );

    \I__622\ : LocalMux
    port map (
            O => \N__4204\,
            I => \uut.pc.G_26_i_a4_5\
        );

    \I__621\ : InMux
    port map (
            O => \N__4201\,
            I => \N__4195\
        );

    \I__620\ : InMux
    port map (
            O => \N__4200\,
            I => \N__4195\
        );

    \I__619\ : LocalMux
    port map (
            O => \N__4195\,
            I => \N__4191\
        );

    \I__618\ : InMux
    port map (
            O => \N__4194\,
            I => \N__4188\
        );

    \I__617\ : Odrv4
    port map (
            O => \N__4191\,
            I => \uut.ir_out_m_c_c_0\
        );

    \I__616\ : LocalMux
    port map (
            O => \N__4188\,
            I => \uut.ir_out_m_c_c_0\
        );

    \I__615\ : InMux
    port map (
            O => \N__4183\,
            I => \N__4180\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__4180\,
            I => \N__4177\
        );

    \I__613\ : Odrv4
    port map (
            O => \N__4177\,
            I => \uut.alu_out_m_0_0\
        );

    \I__612\ : InMux
    port map (
            O => \N__4174\,
            I => \N__4171\
        );

    \I__611\ : LocalMux
    port map (
            O => \N__4171\,
            I => \N__4168\
        );

    \I__610\ : Span4Mux_h
    port map (
            O => \N__4168\,
            I => \N__4165\
        );

    \I__609\ : Odrv4
    port map (
            O => \N__4165\,
            I => \uut.alu_out_m_0\
        );

    \I__608\ : CascadeMux
    port map (
            O => \N__4162\,
            I => \uut.pc.program_counter_4_a1_0_0_1_cascade_\
        );

    \I__607\ : InMux
    port map (
            O => \N__4159\,
            I => \N__4156\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__4156\,
            I => \uut.pc.g2_0\
        );

    \I__605\ : InMux
    port map (
            O => \N__4153\,
            I => \N__4150\
        );

    \I__604\ : LocalMux
    port map (
            O => \N__4150\,
            I => \uut.pc.N_77_0\
        );

    \I__603\ : CascadeMux
    port map (
            O => \N__4147\,
            I => \uut.pc.g1_0_cascade_\
        );

    \I__602\ : InMux
    port map (
            O => \N__4144\,
            I => \N__4139\
        );

    \I__601\ : InMux
    port map (
            O => \N__4143\,
            I => \N__4132\
        );

    \I__600\ : InMux
    port map (
            O => \N__4142\,
            I => \N__4129\
        );

    \I__599\ : LocalMux
    port map (
            O => \N__4139\,
            I => \N__4124\
        );

    \I__598\ : InMux
    port map (
            O => \N__4138\,
            I => \N__4121\
        );

    \I__597\ : InMux
    port map (
            O => \N__4137\,
            I => \N__4118\
        );

    \I__596\ : CascadeMux
    port map (
            O => \N__4136\,
            I => \N__4113\
        );

    \I__595\ : InMux
    port map (
            O => \N__4135\,
            I => \N__4110\
        );

    \I__594\ : LocalMux
    port map (
            O => \N__4132\,
            I => \N__4107\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__4129\,
            I => \N__4104\
        );

    \I__592\ : CascadeMux
    port map (
            O => \N__4128\,
            I => \N__4098\
        );

    \I__591\ : InMux
    port map (
            O => \N__4127\,
            I => \N__4095\
        );

    \I__590\ : Span4Mux_h
    port map (
            O => \N__4124\,
            I => \N__4092\
        );

    \I__589\ : LocalMux
    port map (
            O => \N__4121\,
            I => \N__4087\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__4118\,
            I => \N__4087\
        );

    \I__587\ : InMux
    port map (
            O => \N__4117\,
            I => \N__4080\
        );

    \I__586\ : InMux
    port map (
            O => \N__4116\,
            I => \N__4080\
        );

    \I__585\ : InMux
    port map (
            O => \N__4113\,
            I => \N__4080\
        );

    \I__584\ : LocalMux
    port map (
            O => \N__4110\,
            I => \N__4073\
        );

    \I__583\ : Span4Mux_v
    port map (
            O => \N__4107\,
            I => \N__4073\
        );

    \I__582\ : Span4Mux_v
    port map (
            O => \N__4104\,
            I => \N__4073\
        );

    \I__581\ : InMux
    port map (
            O => \N__4103\,
            I => \N__4070\
        );

    \I__580\ : InMux
    port map (
            O => \N__4102\,
            I => \N__4067\
        );

    \I__579\ : InMux
    port map (
            O => \N__4101\,
            I => \N__4062\
        );

    \I__578\ : InMux
    port map (
            O => \N__4098\,
            I => \N__4062\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__4095\,
            I => \uut.ir_out_7\
        );

    \I__576\ : Odrv4
    port map (
            O => \N__4092\,
            I => \uut.ir_out_7\
        );

    \I__575\ : Odrv12
    port map (
            O => \N__4087\,
            I => \uut.ir_out_7\
        );

    \I__574\ : LocalMux
    port map (
            O => \N__4080\,
            I => \uut.ir_out_7\
        );

    \I__573\ : Odrv4
    port map (
            O => \N__4073\,
            I => \uut.ir_out_7\
        );

    \I__572\ : LocalMux
    port map (
            O => \N__4070\,
            I => \uut.ir_out_7\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__4067\,
            I => \uut.ir_out_7\
        );

    \I__570\ : LocalMux
    port map (
            O => \N__4062\,
            I => \uut.ir_out_7\
        );

    \I__569\ : InMux
    port map (
            O => \N__4045\,
            I => \N__4039\
        );

    \I__568\ : InMux
    port map (
            O => \N__4044\,
            I => \N__4034\
        );

    \I__567\ : InMux
    port map (
            O => \N__4043\,
            I => \N__4034\
        );

    \I__566\ : InMux
    port map (
            O => \N__4042\,
            I => \N__4031\
        );

    \I__565\ : LocalMux
    port map (
            O => \N__4039\,
            I => \N__4028\
        );

    \I__564\ : LocalMux
    port map (
            O => \N__4034\,
            I => \N__4025\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__4031\,
            I => \N__4014\
        );

    \I__562\ : Span4Mux_h
    port map (
            O => \N__4028\,
            I => \N__4014\
        );

    \I__561\ : Span4Mux_v
    port map (
            O => \N__4025\,
            I => \N__4011\
        );

    \I__560\ : InMux
    port map (
            O => \N__4024\,
            I => \N__4006\
        );

    \I__559\ : InMux
    port map (
            O => \N__4023\,
            I => \N__4006\
        );

    \I__558\ : InMux
    port map (
            O => \N__4022\,
            I => \N__4003\
        );

    \I__557\ : InMux
    port map (
            O => \N__4021\,
            I => \N__3996\
        );

    \I__556\ : InMux
    port map (
            O => \N__4020\,
            I => \N__3996\
        );

    \I__555\ : InMux
    port map (
            O => \N__4019\,
            I => \N__3996\
        );

    \I__554\ : Odrv4
    port map (
            O => \N__4014\,
            I => \uut.ir_out_6\
        );

    \I__553\ : Odrv4
    port map (
            O => \N__4011\,
            I => \uut.ir_out_6\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__4006\,
            I => \uut.ir_out_6\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__4003\,
            I => \uut.ir_out_6\
        );

    \I__550\ : LocalMux
    port map (
            O => \N__3996\,
            I => \uut.ir_out_6\
        );

    \I__549\ : InMux
    port map (
            O => \N__3985\,
            I => \N__3982\
        );

    \I__548\ : LocalMux
    port map (
            O => \N__3982\,
            I => \uut.AR_BUF.g0_3_a10_1Z0Z_1\
        );

    \I__547\ : InMux
    port map (
            O => \N__3979\,
            I => \N__3975\
        );

    \I__546\ : InMux
    port map (
            O => \N__3978\,
            I => \N__3972\
        );

    \I__545\ : LocalMux
    port map (
            O => \N__3975\,
            I => \N__3969\
        );

    \I__544\ : LocalMux
    port map (
            O => \N__3972\,
            I => \N__3966\
        );

    \I__543\ : Odrv12
    port map (
            O => \N__3969\,
            I => \uut.D_1_0\
        );

    \I__542\ : Odrv4
    port map (
            O => \N__3966\,
            I => \uut.D_1_0\
        );

    \I__541\ : CascadeMux
    port map (
            O => \N__3961\,
            I => \uut.AR_BUF.g0_3_a10_0Z0Z_2_cascade_\
        );

    \I__540\ : InMux
    port map (
            O => \N__3958\,
            I => \N__3955\
        );

    \I__539\ : LocalMux
    port map (
            O => \N__3955\,
            I => \uut.AR_BUF.g0_3Z0Z_0\
        );

    \I__538\ : CascadeMux
    port map (
            O => \N__3952\,
            I => \uut.ir_out_m_c_d_0_cascade_\
        );

    \I__537\ : InMux
    port map (
            O => \N__3949\,
            I => \N__3946\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__3946\,
            I => \uut.AR_BUF.out_1_2_ivZ0Z_2\
        );

    \I__535\ : CascadeMux
    port map (
            O => \N__3943\,
            I => \N__3940\
        );

    \I__534\ : InMux
    port map (
            O => \N__3940\,
            I => \N__3937\
        );

    \I__533\ : LocalMux
    port map (
            O => \N__3937\,
            I => \N__3934\
        );

    \I__532\ : Odrv4
    port map (
            O => \N__3934\,
            I => \uut.AR_BUF.g0_1_a10_4Z0Z_1\
        );

    \I__531\ : CascadeMux
    port map (
            O => \N__3931\,
            I => \uut.AR_BUF.g0_3Z0Z_2_cascade_\
        );

    \I__530\ : CascadeMux
    port map (
            O => \N__3928\,
            I => \uut.AR_BUF.g0_3Z0Z_6_cascade_\
        );

    \I__529\ : InMux
    port map (
            O => \N__3925\,
            I => \N__3920\
        );

    \I__528\ : InMux
    port map (
            O => \N__3924\,
            I => \N__3915\
        );

    \I__527\ : InMux
    port map (
            O => \N__3923\,
            I => \N__3915\
        );

    \I__526\ : LocalMux
    port map (
            O => \N__3920\,
            I => \uut.AR_out_0\
        );

    \I__525\ : LocalMux
    port map (
            O => \N__3915\,
            I => \uut.AR_out_0\
        );

    \I__524\ : CascadeMux
    port map (
            O => \N__3910\,
            I => \uut.seq.counter.un4_ACC_LD_cascade_\
        );

    \I__523\ : CascadeMux
    port map (
            O => \N__3907\,
            I => \N__3904\
        );

    \I__522\ : InMux
    port map (
            O => \N__3904\,
            I => \N__3901\
        );

    \I__521\ : LocalMux
    port map (
            O => \N__3901\,
            I => \N__3898\
        );

    \I__520\ : Span4Mux_v
    port map (
            O => \N__3898\,
            I => \N__3895\
        );

    \I__519\ : Odrv4
    port map (
            O => \N__3895\,
            I => \uut.seq.counter.ACC_LD_0_0\
        );

    \I__518\ : InMux
    port map (
            O => \N__3892\,
            I => \N__3888\
        );

    \I__517\ : InMux
    port map (
            O => \N__3891\,
            I => \N__3885\
        );

    \I__516\ : LocalMux
    port map (
            O => \N__3888\,
            I => \N__3880\
        );

    \I__515\ : LocalMux
    port map (
            O => \N__3885\,
            I => \N__3877\
        );

    \I__514\ : InMux
    port map (
            O => \N__3884\,
            I => \N__3874\
        );

    \I__513\ : InMux
    port map (
            O => \N__3883\,
            I => \N__3871\
        );

    \I__512\ : Span4Mux_v
    port map (
            O => \N__3880\,
            I => \N__3868\
        );

    \I__511\ : Span4Mux_h
    port map (
            O => \N__3877\,
            I => \N__3863\
        );

    \I__510\ : LocalMux
    port map (
            O => \N__3874\,
            I => \N__3863\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__3871\,
            I => \uut.N_2_0\
        );

    \I__508\ : Odrv4
    port map (
            O => \N__3868\,
            I => \uut.N_2_0\
        );

    \I__507\ : Odrv4
    port map (
            O => \N__3863\,
            I => \uut.N_2_0\
        );

    \I__506\ : InMux
    port map (
            O => \N__3856\,
            I => \N__3850\
        );

    \I__505\ : InMux
    port map (
            O => \N__3855\,
            I => \N__3850\
        );

    \I__504\ : LocalMux
    port map (
            O => \N__3850\,
            I => \N__3844\
        );

    \I__503\ : InMux
    port map (
            O => \N__3849\,
            I => \N__3841\
        );

    \I__502\ : InMux
    port map (
            O => \N__3848\,
            I => \N__3838\
        );

    \I__501\ : InMux
    port map (
            O => \N__3847\,
            I => \N__3835\
        );

    \I__500\ : Odrv4
    port map (
            O => \N__3844\,
            I => \uut.q_ret_1_fast_0\
        );

    \I__499\ : LocalMux
    port map (
            O => \N__3841\,
            I => \uut.q_ret_1_fast_0\
        );

    \I__498\ : LocalMux
    port map (
            O => \N__3838\,
            I => \uut.q_ret_1_fast_0\
        );

    \I__497\ : LocalMux
    port map (
            O => \N__3835\,
            I => \uut.q_ret_1_fast_0\
        );

    \I__496\ : CascadeMux
    port map (
            O => \N__3826\,
            I => \uut.AR_BUF.g0_3Z0Z_3_cascade_\
        );

    \I__495\ : InMux
    port map (
            O => \N__3823\,
            I => \N__3820\
        );

    \I__494\ : LocalMux
    port map (
            O => \N__3820\,
            I => \N__3817\
        );

    \I__493\ : Odrv4
    port map (
            O => \N__3817\,
            I => \uut.AR_BUF.out_1_2_ivZ0Z_1\
        );

    \I__492\ : InMux
    port map (
            O => \N__3814\,
            I => \N__3811\
        );

    \I__491\ : LocalMux
    port map (
            O => \N__3811\,
            I => \N__3807\
        );

    \I__490\ : InMux
    port map (
            O => \N__3810\,
            I => \N__3804\
        );

    \I__489\ : Span4Mux_v
    port map (
            O => \N__3807\,
            I => \N__3798\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__3804\,
            I => \N__3798\
        );

    \I__487\ : CascadeMux
    port map (
            O => \N__3803\,
            I => \N__3794\
        );

    \I__486\ : Span4Mux_v
    port map (
            O => \N__3798\,
            I => \N__3791\
        );

    \I__485\ : InMux
    port map (
            O => \N__3797\,
            I => \N__3788\
        );

    \I__484\ : InMux
    port map (
            O => \N__3794\,
            I => \N__3785\
        );

    \I__483\ : Odrv4
    port map (
            O => \N__3791\,
            I => \uut.un1_HLT_1\
        );

    \I__482\ : LocalMux
    port map (
            O => \N__3788\,
            I => \uut.un1_HLT_1\
        );

    \I__481\ : LocalMux
    port map (
            O => \N__3785\,
            I => \uut.un1_HLT_1\
        );

    \I__480\ : InMux
    port map (
            O => \N__3778\,
            I => \N__3771\
        );

    \I__479\ : InMux
    port map (
            O => \N__3777\,
            I => \N__3771\
        );

    \I__478\ : InMux
    port map (
            O => \N__3776\,
            I => \N__3768\
        );

    \I__477\ : LocalMux
    port map (
            O => \N__3771\,
            I => \N__3765\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__3768\,
            I => \uut.N_5_0\
        );

    \I__475\ : Odrv4
    port map (
            O => \N__3765\,
            I => \uut.N_5_0\
        );

    \I__474\ : InMux
    port map (
            O => \N__3760\,
            I => \N__3757\
        );

    \I__473\ : LocalMux
    port map (
            O => \N__3757\,
            I => \N__3754\
        );

    \I__472\ : Span4Mux_h
    port map (
            O => \N__3754\,
            I => \N__3751\
        );

    \I__471\ : Odrv4
    port map (
            O => \N__3751\,
            I => \uut.bus_6\
        );

    \I__470\ : InMux
    port map (
            O => \N__3748\,
            I => \N__3745\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3745\,
            I => \N__3742\
        );

    \I__468\ : Span4Mux_s2_v
    port map (
            O => \N__3742\,
            I => \N__3739\
        );

    \I__467\ : Odrv4
    port map (
            O => \N__3739\,
            I => \uut.bus_7\
        );

    \I__466\ : CascadeMux
    port map (
            O => \N__3736\,
            I => \uut.seq.D_2_0_x_cascade_\
        );

    \I__465\ : CascadeMux
    port map (
            O => \N__3733\,
            I => \N__3728\
        );

    \I__464\ : CascadeMux
    port map (
            O => \N__3732\,
            I => \N__3725\
        );

    \I__463\ : InMux
    port map (
            O => \N__3731\,
            I => \N__3722\
        );

    \I__462\ : InMux
    port map (
            O => \N__3728\,
            I => \N__3719\
        );

    \I__461\ : InMux
    port map (
            O => \N__3725\,
            I => \N__3716\
        );

    \I__460\ : LocalMux
    port map (
            O => \N__3722\,
            I => \uut.q_0_fast\
        );

    \I__459\ : LocalMux
    port map (
            O => \N__3719\,
            I => \uut.q_0_fast\
        );

    \I__458\ : LocalMux
    port map (
            O => \N__3716\,
            I => \uut.q_0_fast\
        );

    \I__457\ : InMux
    port map (
            O => \N__3709\,
            I => \N__3703\
        );

    \I__456\ : InMux
    port map (
            O => \N__3708\,
            I => \N__3703\
        );

    \I__455\ : LocalMux
    port map (
            O => \N__3703\,
            I => \N__3700\
        );

    \I__454\ : Odrv4
    port map (
            O => \N__3700\,
            I => \uut.data_1_2_ivdup\
        );

    \I__453\ : CascadeMux
    port map (
            O => \N__3697\,
            I => \uut.IR.ir_out_m_c_d_1_3_cascade_\
        );

    \I__452\ : CascadeMux
    port map (
            O => \N__3694\,
            I => \uut.ir_out_m_c_d_3_cascade_\
        );

    \I__451\ : InMux
    port map (
            O => \N__3691\,
            I => \N__3688\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__3688\,
            I => \uut.seq.counter.T_2_rep1_RNIGC8CZ0Z1\
        );

    \I__449\ : CascadeMux
    port map (
            O => \N__3685\,
            I => \uut.seq.un13_ACC_LD_xZ0Z1_cascade_\
        );

    \I__448\ : CascadeMux
    port map (
            O => \N__3682\,
            I => \uut.seq.counter.T_2_rep1_RNI8TEZ0Z81_cascade_\
        );

    \I__447\ : CascadeMux
    port map (
            O => \N__3679\,
            I => \uut.seq.counter.un2_MAR_LD_cascade_\
        );

    \I__446\ : CascadeMux
    port map (
            O => \N__3676\,
            I => \uut.D_1_0_cascade_\
        );

    \I__445\ : InMux
    port map (
            O => \N__3673\,
            I => \N__3670\
        );

    \I__444\ : LocalMux
    port map (
            O => \N__3670\,
            I => \uut.seq.q_ret_RNI52E81Z0Z_0\
        );

    \I__443\ : CascadeMux
    port map (
            O => \N__3667\,
            I => \uut.T_2_rep1_RNI6BLF1_cascade_\
        );

    \I__442\ : CascadeMux
    port map (
            O => \N__3664\,
            I => \N__3661\
        );

    \I__441\ : InMux
    port map (
            O => \N__3661\,
            I => \N__3658\
        );

    \I__440\ : LocalMux
    port map (
            O => \N__3658\,
            I => \N__3655\
        );

    \I__439\ : Span4Mux_h
    port map (
            O => \N__3655\,
            I => \N__3652\
        );

    \I__438\ : Odrv4
    port map (
            O => \N__3652\,
            I => \uut.un17_IR_OE_0\
        );

    \I__437\ : InMux
    port map (
            O => \N__3649\,
            I => \N__3645\
        );

    \I__436\ : CascadeMux
    port map (
            O => \N__3648\,
            I => \N__3642\
        );

    \I__435\ : LocalMux
    port map (
            O => \N__3645\,
            I => \N__3639\
        );

    \I__434\ : InMux
    port map (
            O => \N__3642\,
            I => \N__3636\
        );

    \I__433\ : Odrv4
    port map (
            O => \N__3639\,
            I => \uut.ir_out_m_d_0\
        );

    \I__432\ : LocalMux
    port map (
            O => \N__3636\,
            I => \uut.ir_out_m_d_0\
        );

    \I__431\ : CascadeMux
    port map (
            O => \N__3631\,
            I => \uut.pc.N_4_i_1_cascade_\
        );

    \I__430\ : InMux
    port map (
            O => \N__3628\,
            I => \N__3624\
        );

    \I__429\ : InMux
    port map (
            O => \N__3627\,
            I => \N__3621\
        );

    \I__428\ : LocalMux
    port map (
            O => \N__3624\,
            I => \uut.alu_out_m_2\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__3621\,
            I => \uut.alu_out_m_2\
        );

    \I__426\ : CascadeMux
    port map (
            O => \N__3616\,
            I => \uut.ALU_main.N_43_0_cascade_\
        );

    \I__425\ : CascadeMux
    port map (
            O => \N__3613\,
            I => \uut.T_1_fast_RNIVM0N3_0_cascade_\
        );

    \I__424\ : InMux
    port map (
            O => \N__3610\,
            I => \N__3607\
        );

    \I__423\ : LocalMux
    port map (
            O => \N__3607\,
            I => \uut.pc.N_11\
        );

    \I__422\ : CascadeMux
    port map (
            O => \N__3604\,
            I => \uut.AR_BUF.N_13_cascade_\
        );

    \I__421\ : CascadeMux
    port map (
            O => \N__3601\,
            I => \uut.AR_BUF.g0_1_0Z0Z_5_cascade_\
        );

    \I__420\ : InMux
    port map (
            O => \N__3598\,
            I => \N__3595\
        );

    \I__419\ : LocalMux
    port map (
            O => \N__3595\,
            I => \uut.AR_BUF.g0_1_0Z0Z_1\
        );

    \I__418\ : CascadeMux
    port map (
            O => \N__3592\,
            I => \N__3589\
        );

    \I__417\ : InMux
    port map (
            O => \N__3589\,
            I => \N__3585\
        );

    \I__416\ : CascadeMux
    port map (
            O => \N__3588\,
            I => \N__3581\
        );

    \I__415\ : LocalMux
    port map (
            O => \N__3585\,
            I => \N__3578\
        );

    \I__414\ : InMux
    port map (
            O => \N__3584\,
            I => \N__3573\
        );

    \I__413\ : InMux
    port map (
            O => \N__3581\,
            I => \N__3573\
        );

    \I__412\ : Span4Mux_v
    port map (
            O => \N__3578\,
            I => \N__3570\
        );

    \I__411\ : LocalMux
    port map (
            O => \N__3573\,
            I => \uut.AR_out_1\
        );

    \I__410\ : Odrv4
    port map (
            O => \N__3570\,
            I => \uut.AR_out_1\
        );

    \I__409\ : InMux
    port map (
            O => \N__3565\,
            I => \N__3562\
        );

    \I__408\ : LocalMux
    port map (
            O => \N__3562\,
            I => \uut.AR_BUF.g0_1_0_4_0\
        );

    \I__407\ : CascadeMux
    port map (
            O => \N__3559\,
            I => \N__3554\
        );

    \I__406\ : CascadeMux
    port map (
            O => \N__3558\,
            I => \N__3548\
        );

    \I__405\ : InMux
    port map (
            O => \N__3557\,
            I => \N__3545\
        );

    \I__404\ : InMux
    port map (
            O => \N__3554\,
            I => \N__3541\
        );

    \I__403\ : InMux
    port map (
            O => \N__3553\,
            I => \N__3534\
        );

    \I__402\ : InMux
    port map (
            O => \N__3552\,
            I => \N__3534\
        );

    \I__401\ : InMux
    port map (
            O => \N__3551\,
            I => \N__3534\
        );

    \I__400\ : InMux
    port map (
            O => \N__3548\,
            I => \N__3531\
        );

    \I__399\ : LocalMux
    port map (
            O => \N__3545\,
            I => \N__3528\
        );

    \I__398\ : InMux
    port map (
            O => \N__3544\,
            I => \N__3525\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__3541\,
            I => \N__3522\
        );

    \I__396\ : LocalMux
    port map (
            O => \N__3534\,
            I => \N__3517\
        );

    \I__395\ : LocalMux
    port map (
            O => \N__3531\,
            I => \N__3517\
        );

    \I__394\ : Sp12to4
    port map (
            O => \N__3528\,
            I => \N__3512\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__3525\,
            I => \N__3512\
        );

    \I__392\ : Span4Mux_v
    port map (
            O => \N__3522\,
            I => \N__3507\
        );

    \I__391\ : Span4Mux_v
    port map (
            O => \N__3517\,
            I => \N__3507\
        );

    \I__390\ : Odrv12
    port map (
            O => \N__3512\,
            I => \uut.ir_out_1\
        );

    \I__389\ : Odrv4
    port map (
            O => \N__3507\,
            I => \uut.ir_out_1\
        );

    \I__388\ : InMux
    port map (
            O => \N__3502\,
            I => \N__3499\
        );

    \I__387\ : LocalMux
    port map (
            O => \N__3499\,
            I => \uut.AR_BUF.N_10\
        );

    \I__386\ : InMux
    port map (
            O => \N__3496\,
            I => \N__3493\
        );

    \I__385\ : LocalMux
    port map (
            O => \N__3493\,
            I => \uut.AR_BUF.g0_1_0_0_0\
        );

    \I__384\ : InMux
    port map (
            O => \N__3490\,
            I => \N__3487\
        );

    \I__383\ : LocalMux
    port map (
            O => \N__3487\,
            I => \N__3484\
        );

    \I__382\ : Odrv4
    port map (
            O => \N__3484\,
            I => \uut.AR_BUF.out_1_0_iv_2_1Z0Z_1\
        );

    \I__381\ : CascadeMux
    port map (
            O => \N__3481\,
            I => \uut.AR_BUF.g0_0_a5_0Z0Z_2_cascade_\
        );

    \I__380\ : InMux
    port map (
            O => \N__3478\,
            I => \N__3475\
        );

    \I__379\ : LocalMux
    port map (
            O => \N__3475\,
            I => \N__3472\
        );

    \I__378\ : Odrv12
    port map (
            O => \N__3472\,
            I => \uut.AR_BUF.N_9\
        );

    \I__377\ : CascadeMux
    port map (
            O => \N__3469\,
            I => \N__3466\
        );

    \I__376\ : InMux
    port map (
            O => \N__3466\,
            I => \N__3463\
        );

    \I__375\ : LocalMux
    port map (
            O => \N__3463\,
            I => \uut.AR_BUF.g0_1_a10_3Z0Z_2\
        );

    \I__374\ : InMux
    port map (
            O => \N__3460\,
            I => \N__3457\
        );

    \I__373\ : LocalMux
    port map (
            O => \N__3457\,
            I => \uut.AR_BUF.g0_0_o5_0Z0Z_0\
        );

    \I__372\ : CascadeMux
    port map (
            O => \N__3454\,
            I => \uut.AR_BUF.g0_1_a10_3_cascade_\
        );

    \I__371\ : InMux
    port map (
            O => \N__3451\,
            I => \N__3448\
        );

    \I__370\ : LocalMux
    port map (
            O => \N__3448\,
            I => \uut.AR_BUF.N_7\
        );

    \I__369\ : InMux
    port map (
            O => \N__3445\,
            I => \N__3439\
        );

    \I__368\ : InMux
    port map (
            O => \N__3444\,
            I => \N__3439\
        );

    \I__367\ : LocalMux
    port map (
            O => \N__3439\,
            I => \uut.b_reg_out_4\
        );

    \I__366\ : InMux
    port map (
            O => \N__3436\,
            I => \N__3433\
        );

    \I__365\ : LocalMux
    port map (
            O => \N__3433\,
            I => \N__3430\
        );

    \I__364\ : Odrv12
    port map (
            O => \N__3430\,
            I => \uut.AR_BUF.out_1_0_iv_2Z0Z_0\
        );

    \I__363\ : CascadeMux
    port map (
            O => \N__3427\,
            I => \uut.ir_out_m_d_2_cascade_\
        );

    \I__362\ : CascadeMux
    port map (
            O => \N__3424\,
            I => \N__3421\
        );

    \I__361\ : InMux
    port map (
            O => \N__3421\,
            I => \N__3418\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__3418\,
            I => \uut.ALU_main.N_48\
        );

    \I__359\ : CascadeMux
    port map (
            O => \N__3415\,
            I => \uut.bus_6_cascade_\
        );

    \I__358\ : CascadeMux
    port map (
            O => \N__3412\,
            I => \uut.q_RNIDGA71_cascade_\
        );

    \I__357\ : CascadeMux
    port map (
            O => \N__3409\,
            I => \uut.ALU_main.N_45_cascade_\
        );

    \I__356\ : CascadeMux
    port map (
            O => \N__3406\,
            I => \uut.alu_out_m_4_cascade_\
        );

    \I__355\ : CascadeMux
    port map (
            O => \N__3403\,
            I => \uut.data_1_2_ivdup_cascade_\
        );

    \I__354\ : InMux
    port map (
            O => \N__3400\,
            I => \N__3397\
        );

    \I__353\ : LocalMux
    port map (
            O => \N__3397\,
            I => \uut.N_4_0\
        );

    \I__352\ : InMux
    port map (
            O => \N__3394\,
            I => \N__3391\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__3391\,
            I => \N__3388\
        );

    \I__350\ : Span4Mux_h
    port map (
            O => \N__3388\,
            I => \N__3385\
        );

    \I__349\ : Odrv4
    port map (
            O => \N__3385\,
            I => \uut.data_1_2_iv_0\
        );

    \I__348\ : CascadeMux
    port map (
            O => \N__3382\,
            I => \uut.program_counter_m_2_cascade_\
        );

    \I__347\ : InMux
    port map (
            O => \N__3379\,
            I => \N__3376\
        );

    \I__346\ : LocalMux
    port map (
            O => \N__3376\,
            I => \uut.AR_BUF.N_8\
        );

    \I__345\ : CascadeMux
    port map (
            O => \N__3373\,
            I => \N__3370\
        );

    \I__344\ : InMux
    port map (
            O => \N__3370\,
            I => \N__3367\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__3367\,
            I => \uut.program_counter_m_2\
        );

    \I__342\ : InMux
    port map (
            O => \N__3364\,
            I => \N__3361\
        );

    \I__341\ : LocalMux
    port map (
            O => \N__3361\,
            I => \uut.AR_BUF.g0_0_0Z0Z_1\
        );

    \I__340\ : CascadeMux
    port map (
            O => \N__3358\,
            I => \uut.out_1_0_ivdup_2_cascade_\
        );

    \I__339\ : InMux
    port map (
            O => \N__3355\,
            I => \N__3352\
        );

    \I__338\ : LocalMux
    port map (
            O => \N__3352\,
            I => \uut.ALU_main.N_43\
        );

    \I__337\ : InMux
    port map (
            O => \N__3349\,
            I => \N__3346\
        );

    \I__336\ : LocalMux
    port map (
            O => \N__3346\,
            I => \uut.ir_out_m_d_1\
        );

    \I__335\ : CascadeMux
    port map (
            O => \N__3343\,
            I => \uut.acc_out_m_7_cascade_\
        );

    \I__334\ : CascadeMux
    port map (
            O => \N__3340\,
            I => \uut.bus_7_cascade_\
        );

    \I__333\ : InMux
    port map (
            O => \N__3337\,
            I => \N__3334\
        );

    \I__332\ : LocalMux
    port map (
            O => \N__3334\,
            I => \N__3331\
        );

    \I__331\ : Odrv4
    port map (
            O => \N__3331\,
            I => \uut.N_1_0\
        );

    \I__330\ : IoInMux
    port map (
            O => \N__3328\,
            I => \N__3325\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__3325\,
            I => \N__3322\
        );

    \I__328\ : Span4Mux_s2_h
    port map (
            O => \N__3322\,
            I => \N__3319\
        );

    \I__327\ : Span4Mux_v
    port map (
            O => \N__3319\,
            I => \N__3315\
        );

    \I__326\ : CascadeMux
    port map (
            O => \N__3318\,
            I => \N__3312\
        );

    \I__325\ : Span4Mux_h
    port map (
            O => \N__3315\,
            I => \N__3309\
        );

    \I__324\ : InMux
    port map (
            O => \N__3312\,
            I => \N__3306\
        );

    \I__323\ : Odrv4
    port map (
            O => \N__3309\,
            I => \LED5_c\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__3306\,
            I => \LED5_c\
        );

    \I__321\ : CascadeMux
    port map (
            O => \N__3301\,
            I => \uut.out_1_2_iv_3_cascade_\
        );

    \I__320\ : IoInMux
    port map (
            O => \N__3298\,
            I => \N__3295\
        );

    \I__319\ : LocalMux
    port map (
            O => \N__3295\,
            I => \N__3292\
        );

    \I__318\ : Span4Mux_s2_h
    port map (
            O => \N__3292\,
            I => \N__3289\
        );

    \I__317\ : Span4Mux_v
    port map (
            O => \N__3289\,
            I => \N__3285\
        );

    \I__316\ : InMux
    port map (
            O => \N__3288\,
            I => \N__3282\
        );

    \I__315\ : Odrv4
    port map (
            O => \N__3285\,
            I => \LED1_c\
        );

    \I__314\ : LocalMux
    port map (
            O => \N__3282\,
            I => \LED1_c\
        );

    \I__313\ : CascadeMux
    port map (
            O => \N__3277\,
            I => \uut.ALU_main.N_47_cascade_\
        );

    \I__312\ : CascadeMux
    port map (
            O => \N__3274\,
            I => \uut.seq.un1_HLT_1_reti_cascade_\
        );

    \I__311\ : InMux
    port map (
            O => \N__3271\,
            I => \N__3268\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__3268\,
            I => \N__3265\
        );

    \I__309\ : Odrv4
    port map (
            O => \N__3265\,
            I => \uut.un1_HLT_0\
        );

    \I__308\ : CascadeMux
    port map (
            O => \N__3262\,
            I => \uut.ALU_main.N_46_cascade_\
        );

    \I__307\ : CascadeMux
    port map (
            O => \N__3259\,
            I => \uut.alu_out_m_5_cascade_\
        );

    \I__306\ : CascadeMux
    port map (
            O => \N__3256\,
            I => \uut.bus_5_cascade_\
        );

    \I__305\ : CascadeMux
    port map (
            O => \N__3253\,
            I => \uut.alu_out_m_7_cascade_\
        );

    \I__304\ : CascadeMux
    port map (
            O => \N__3250\,
            I => \uut.AR_BUF.out_1_1_iv_3_1Z0Z_0_cascade_\
        );

    \I__303\ : CascadeMux
    port map (
            O => \N__3247\,
            I => \uut.AR_BUF.out_1_1_ivZ0Z_0_cascade_\
        );

    \I__302\ : CascadeMux
    port map (
            O => \N__3244\,
            I => \uut.out_1_1_iv_2_cascade_\
        );

    \I__301\ : InMux
    port map (
            O => \N__3241\,
            I => \N__3238\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__3238\,
            I => \G_138\
        );

    \I__299\ : CascadeMux
    port map (
            O => \N__3235\,
            I => \G_138_cascade_\
        );

    \I__298\ : IoInMux
    port map (
            O => \N__3232\,
            I => \N__3229\
        );

    \I__297\ : LocalMux
    port map (
            O => \N__3229\,
            I => \N__3226\
        );

    \I__296\ : Odrv12
    port map (
            O => \N__3226\,
            I => \uut.buf_clk_1\
        );

    \INVuut.mar.ff4.q_neC\ : INV
    port map (
            O => \INVuut.mar.ff4.q_neC_net\,
            I => \N__5658\
        );

    \INVuut.out_reg.ff4.qC\ : INV
    port map (
            O => \INVuut.out_reg.ff4.qC_net\,
            I => \N__5656\
        );

    \INVuut.seq.counter.T_1_0C\ : INV
    port map (
            O => \INVuut.seq.counter.T_1_0C_net\,
            I => \N__5652\
        );

    \INVuut.AR.ff4.q_neC\ : INV
    port map (
            O => \INVuut.AR.ff4.q_neC_net\,
            I => \N__5649\
        );

    \INVuut.AR.ff3.qC\ : INV
    port map (
            O => \INVuut.AR.ff3.qC_net\,
            I => \N__5645\
        );

    \INVuut.IR.ff3.qC\ : INV
    port map (
            O => \INVuut.IR.ff3.qC_net\,
            I => \N__5659\
        );

    \INVuut.b_reg.ff1.qC\ : INV
    port map (
            O => \INVuut.b_reg.ff1.qC_net\,
            I => \N__5657\
        );

    \INVuut.out_reg.ff3.qC\ : INV
    port map (
            O => \INVuut.out_reg.ff3.qC_net\,
            I => \N__5655\
        );

    \INVuut.acc.ff4.qC\ : INV
    port map (
            O => \INVuut.acc.ff4.qC_net\,
            I => \N__5651\
        );

    \INVuut.mar.ff2.q_neC\ : INV
    port map (
            O => \INVuut.mar.ff2.q_neC_net\,
            I => \N__5644\
        );

    \INVuut.seq.counter.T_1_1C\ : INV
    port map (
            O => \INVuut.seq.counter.T_1_1C_net\,
            I => \N__5641\
        );

    \INVuut.seq.counter.T_1_4C\ : INV
    port map (
            O => \INVuut.seq.counter.T_1_4C_net\,
            I => \N__5637\
        );

    \INVuut.IR.ff6.q_0_fastC\ : INV
    port map (
            O => \INVuut.IR.ff6.q_0_fastC_net\,
            I => \N__5654\
        );

    \INVuut.b_reg.ff4.qC\ : INV
    port map (
            O => \INVuut.b_reg.ff4.qC_net\,
            I => \N__5640\
        );

    \INVuut.AR.ff1.q_neC\ : INV
    port map (
            O => \INVuut.AR.ff1.q_neC_net\,
            I => \N__5635\
        );

    \INVuut.acc.ff1.qC\ : INV
    port map (
            O => \INVuut.acc.ff1.qC_net\,
            I => \N__5636\
        );

    \INVuut.seq.counter.T_1_fast_3C\ : INV
    port map (
            O => \INVuut.seq.counter.T_1_fast_3C_net\,
            I => \N__5653\
        );

    \INVuut.IR.ff5.q_0_rep1C\ : INV
    port map (
            O => \INVuut.IR.ff5.q_0_rep1C_net\,
            I => \N__5650\
        );

    \INVuut.IR.ff7.q_ret_1_fastC\ : INV
    port map (
            O => \INVuut.IR.ff7.q_ret_1_fastC_net\,
            I => \N__5647\
        );

    \INVuut.IR.ff4.q_neC\ : INV
    port map (
            O => \INVuut.IR.ff4.q_neC_net\,
            I => \N__5643\
        );

    \INVuut.b_reg.ff3.qC\ : INV
    port map (
            O => \INVuut.b_reg.ff3.qC_net\,
            I => \N__5634\
        );

    \INVuut.IR.ff1.q_neC\ : INV
    port map (
            O => \INVuut.IR.ff1.q_neC_net\,
            I => \N__5646\
        );

    \INVuut.seq.q_retC\ : INV
    port map (
            O => \INVuut.seq.q_retC_net\,
            I => \N__5642\
        );

    \INVuut.IR.ff5.q_0_neC\ : INV
    port map (
            O => \INVuut.IR.ff5.q_0_neC_net\,
            I => \N__5639\
        );

    \INVuut.b_reg.ff5.qC\ : INV
    port map (
            O => \INVuut.b_reg.ff5.qC_net\,
            I => \N__5633\
        );

    \INVuut.acc.ff3.qC\ : INV
    port map (
            O => \INVuut.acc.ff3.qC_net\,
            I => \N__5624\
        );

    \INVuut.out_reg.ff1.qC\ : INV
    port map (
            O => \INVuut.out_reg.ff1.qC_net\,
            I => \N__5628\
        );

    \INVuut.out_reg.ff5.qC\ : INV
    port map (
            O => \INVuut.out_reg.ff5.qC_net\,
            I => \N__5638\
        );

    \INVuut.b_reg.ff8.qC\ : INV
    port map (
            O => \INVuut.b_reg.ff8.qC_net\,
            I => \N__5632\
        );

    \INVuut.seq.q_ret_1C\ : INV
    port map (
            O => \INVuut.seq.q_ret_1C_net\,
            I => \N__5630\
        );

    \INVuut.AR.ff2.qC\ : INV
    port map (
            O => \INVuut.AR.ff2.qC_net\,
            I => \N__5625\
        );

    \INVuut.acc.ff2.qC\ : INV
    port map (
            O => \INVuut.acc.ff2.qC_net\,
            I => \N__5623\
        );

    \INVuut.b_reg.ff7.qC\ : INV
    port map (
            O => \INVuut.b_reg.ff7.qC_net\,
            I => \N__5629\
        );

    \INVuut.b_reg.ff6.qC\ : INV
    port map (
            O => \INVuut.b_reg.ff6.qC_net\,
            I => \N__5626\
        );

    \IN_MUX_bfv_9_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_9_12_0_\
        );

    \IN_MUX_bfv_9_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \uut.ALU_main.un1_A_cry_6\,
            carryinitout => \bfn_9_13_0_\
        );

    \uut.buf_clk_1_inferred_clock_0_RNIQBSF\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__3232\,
            GLOBALBUFFEROUTPUT => \uut.buf_clk_1_g\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \N_62_i_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3241\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \G_138\,
            ltout => \G_138_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.buf_clk_1_inferred_clock_0_RNO_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000001010000"
        )
    port map (
            in0 => \N__3271\,
            in1 => \_gnd_net_\,
            in2 => \N__3235\,
            in3 => \_gnd_net_\,
            lcout => \uut.buf_clk_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.b_reg.ff6.q_LC_5_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__6101\,
            in1 => \N__6128\,
            in2 => \N__6079\,
            in3 => \N__9044\,
            lcout => \uut.b_reg_out_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.b_reg.ff6.qC_net\,
            ce => \N__7515\,
            sr => \_gnd_net_\
        );

    \uut.b_reg.ff7.q_LC_5_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__6363\,
            in1 => \N__6402\,
            in2 => \N__6331\,
            in3 => \N__9045\,
            lcout => \uut.b_reg_out_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.b_reg.ff7.qC_net\,
            ce => \N__7514\,
            sr => \_gnd_net_\
        );

    \uut.acc.ff2.q_LC_6_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7684\,
            in1 => \N__7644\,
            in2 => \_gnd_net_\,
            in3 => \N__7579\,
            lcout => \uut.acc_out_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.acc.ff2.qC_net\,
            ce => \N__5833\,
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.out_1_1_iv_3_1_0_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__5171\,
            in1 => \N__8282\,
            in2 => \N__3588\,
            in3 => \N__7783\,
            lcout => OPEN,
            ltout => \uut.AR_BUF.out_1_1_iv_3_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.out_1_1_iv_0_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101111111010"
        )
    port map (
            in0 => \N__5750\,
            in1 => \N__7102\,
            in2 => \N__3250\,
            in3 => \N__3557\,
            lcout => OPEN,
            ltout => \uut.AR_BUF.out_1_1_ivZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.out_1_1_iv_2_LC_6_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110001"
        )
    port map (
            in0 => \N__9072\,
            in1 => \N__6817\,
            in2 => \N__3247\,
            in3 => \N__3349\,
            lcout => OPEN,
            ltout => \uut.out_1_1_iv_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR.ff2.q_LC_6_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101111001000"
        )
    port map (
            in0 => \N__7692\,
            in1 => \N__8032\,
            in2 => \N__3244\,
            in3 => \N__3584\,
            lcout => \uut.AR_out_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.AR.ff2.qC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.acc.ff6.q_RNIEIB71_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6030\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8281\,
            lcout => \uut.acc_out_m_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.ALU_Out_0_6_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001100110"
        )
    port map (
            in0 => \N__6272\,
            in1 => \N__4582\,
            in2 => \_gnd_net_\,
            in3 => \N__6774\,
            lcout => OPEN,
            ltout => \uut.ALU_main.N_47_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_cry_5_c_RNISM3EE_LC_6_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__4615\,
            in1 => \N__6616\,
            in2 => \N__3277\,
            in3 => \N__6492\,
            lcout => \uut.alu_out_m_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_RNIT9ANK_1_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7414\,
            in2 => \_gnd_net_\,
            in3 => \N__3883\,
            lcout => OPEN,
            ltout => \uut.seq.un1_HLT_1_reti_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.q_ret_1_LC_6_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__3776\,
            in1 => \N__3400\,
            in2 => \N__3274\,
            in3 => \N__3337\,
            lcout => \uut.un1_HLT_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.seq.q_ret_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.ALU_Out_0_5_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001100110"
        )
    port map (
            in0 => \N__4554\,
            in1 => \N__6029\,
            in2 => \_gnd_net_\,
            in3 => \N__6766\,
            lcout => OPEN,
            ltout => \uut.ALU_main.N_46_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_cry_4_c_RNIMATDE_LC_6_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__4252\,
            in1 => \N__6620\,
            in2 => \N__3262\,
            in3 => \N__6502\,
            lcout => \uut.alu_out_m_5\,
            ltout => \uut.alu_out_m_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mem.data_1_1_iv_LC_6_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111101"
        )
    port map (
            in0 => \N__6074\,
            in1 => \N__6100\,
            in2 => \N__3259\,
            in3 => \N__9038\,
            lcout => \uut.bus_5\,
            ltout => \uut.bus_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff6.q_0_ne_RNIV8OLK_LC_6_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7413\,
            in2 => \N__3256\,
            in3 => \N__4936\,
            lcout => \uut.N_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_cry_6_c_RNIUOL0E_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__4597\,
            in1 => \N__6619\,
            in2 => \N__3424\,
            in3 => \N__6501\,
            lcout => \uut.alu_out_m_7\,
            ltout => \uut.alu_out_m_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.b_reg.ff8.q_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011111011"
        )
    port map (
            in0 => \N__6215\,
            in1 => \N__6889\,
            in2 => \N__3253\,
            in3 => \N__9074\,
            lcout => \uut.b_reg_out_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.b_reg.ff8.qC_net\,
            ce => \N__7503\,
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_RNI5ENL7_3_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__6760\,
            in1 => \N__4768\,
            in2 => \N__3907\,
            in3 => \N__4423\,
            lcout => \uut.ACC_LD_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.acc.ff8.q_RNIGMD71_LC_6_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__6178\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8273\,
            lcout => \uut.acc_out_m_7\,
            ltout => \uut.acc_out_m_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mem.data_1_iv_LC_6_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111101"
        )
    port map (
            in0 => \N__9005\,
            in1 => \N__6194\,
            in2 => \N__3343\,
            in3 => \N__6874\,
            lcout => \uut.bus_7\,
            ltout => \uut.bus_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff8.q_0_ne_RNIB9TFK_LC_6_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4127\,
            in2 => \N__3340\,
            in3 => \N__7415\,
            lcout => \uut.N_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.out_reg.ff5.q_LC_6_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011011000"
        )
    port map (
            in0 => \N__8274\,
            in1 => \N__3394\,
            in2 => \N__3318\,
            in3 => \N__5913\,
            lcout => \LED5_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.out_reg.ff5.qC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_1_a10_3_2_LC_7_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__4701\,
            in1 => \N__3544\,
            in2 => \_gnd_net_\,
            in3 => \N__4137\,
            lcout => \uut.AR_BUF.g0_1_a10_3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.out_1_2_iv_3_LC_7_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__4174\,
            in1 => \N__3823\,
            in2 => \_gnd_net_\,
            in3 => \N__3649\,
            lcout => OPEN,
            ltout => \uut.out_1_2_iv_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.out_reg.ff1.q_LC_7_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011100010"
        )
    port map (
            in0 => \N__3288\,
            in1 => \N__8287\,
            in2 => \N__3301\,
            in3 => \N__9262\,
            lcout => \LED1_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.out_reg.ff1.qC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.acc.ff3.q_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__8098\,
            in1 => \N__3627\,
            in2 => \N__5452\,
            in3 => \N__9073\,
            lcout => \uut.acc_out_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.acc.ff3.qC_net\,
            ce => \N__5845\,
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_0_0_1_LC_7_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__7762\,
            in1 => \N__4466\,
            in2 => \N__7171\,
            in3 => \N__8260\,
            lcout => \uut.AR_BUF.g0_0_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_0_a5_LC_7_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011100000"
        )
    port map (
            in0 => \N__7974\,
            in1 => \N__3460\,
            in2 => \N__7258\,
            in3 => \N__8385\,
            lcout => \uut.AR_BUF.N_8\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_RNIEETC1_0_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__8756\,
            in1 => \N__8659\,
            in2 => \N__5792\,
            in3 => \N__8579\,
            lcout => \uut.program_counter_m_2\,
            ltout => \uut.program_counter_m_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.out_1_0_iv_2_0_LC_7_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7167\,
            in2 => \N__3382\,
            in3 => \N__7764\,
            lcout => \uut.AR_BUF.out_1_0_iv_2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_cry_1_c_RNI46ADE_0_LC_7_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__6618\,
            in1 => \N__3355\,
            in2 => \N__6496\,
            in3 => \N__4303\,
            lcout => \uut.alu_out_m_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_0_0_LC_7_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3379\,
            in1 => \N__3478\,
            in2 => \N__3373\,
            in3 => \N__3364\,
            lcout => \uut.out_1_0_ivdup_2\,
            ltout => \uut.out_1_0_ivdup_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.pc.program_counter_2_LC_7_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110111001"
        )
    port map (
            in0 => \N__5485\,
            in1 => \N__5461\,
            in2 => \N__3358\,
            in3 => \N__7185\,
            lcout => \uut.program_counter_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5627\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.ALU_Out_0_2_LC_7_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001100110"
        )
    port map (
            in0 => \N__4468\,
            in1 => \N__4500\,
            in2 => \_gnd_net_\,
            in3 => \N__6775\,
            lcout => \uut.ALU_main.N_43\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff1.q_ne_RNI2QSE5_LC_7_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100011001100"
        )
    port map (
            in0 => \N__7933\,
            in1 => \N__5302\,
            in2 => \N__7975\,
            in3 => \N__7872\,
            lcout => \uut.ir_out_m_d_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff2.q_ne_RNI3V695_LC_7_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011010000"
        )
    port map (
            in0 => \N__7873\,
            in1 => \N__7934\,
            in2 => \N__3559\,
            in3 => \N__7965\,
            lcout => \uut.ir_out_m_d_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mem.data_1_0_iv_LC_7_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__6395\,
            in1 => \N__6349\,
            in2 => \N__6316\,
            in3 => \N__9046\,
            lcout => \uut.bus_6\,
            ltout => \uut.bus_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff7.q_0_ne_RNI7UKPK_LC_7_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7403\,
            in2 => \N__3415\,
            in3 => \N__4042\,
            lcout => \uut.N_5_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.acc.ff5.q_RNIDGA71_LC_7_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5878\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8271\,
            lcout => \uut.q_RNIDGA71\,
            ltout => \uut.q_RNIDGA71_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.b_reg.ff5.q_LC_7_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110001"
        )
    port map (
            in0 => \N__5948\,
            in1 => \N__9043\,
            in2 => \N__3412\,
            in3 => \N__5905\,
            lcout => \uut.b_reg_out_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.b_reg.ff5.qC_net\,
            ce => \N__7510\,
            sr => \_gnd_net_\
        );

    \uut.ALU_main.ALU_Out_0_4_LC_7_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001100110"
        )
    port map (
            in0 => \N__5877\,
            in1 => \N__3445\,
            in2 => \_gnd_net_\,
            in3 => \N__6767\,
            lcout => OPEN,
            ltout => \uut.ALU_main.N_45_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_cry_3_c_RNIGUMDE_LC_7_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__4264\,
            in1 => \N__6621\,
            in2 => \N__3409\,
            in3 => \N__6475\,
            lcout => \uut.alu_out_m_4\,
            ltout => \uut.alu_out_m_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mem.data_1_2_ivdup_LC_7_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110001"
        )
    port map (
            in0 => \N__9042\,
            in1 => \N__5947\,
            in2 => \N__3406\,
            in3 => \N__5966\,
            lcout => \uut.data_1_2_ivdup\,
            ltout => \uut.data_1_2_ivdup_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff5.q_0_ne_RNINJRHK_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \N__4700\,
            in1 => \_gnd_net_\,
            in2 => \N__3403\,
            in3 => \N__7412\,
            lcout => \uut.N_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mem.data_1_2_iv_0_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010101111"
        )
    port map (
            in0 => \N__5879\,
            in1 => \_gnd_net_\,
            in2 => \N__9071\,
            in3 => \N__5946\,
            lcout => \uut.data_1_2_iv_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_axb_4_l_ofx_LC_7_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100110"
        )
    port map (
            in0 => \N__3444\,
            in1 => \N__4767\,
            in2 => \N__5884\,
            in3 => \N__4419\,
            lcout => \uut.ALU_main.un1_A_axb_4_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff5.q_0_ne_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011111101"
        )
    port map (
            in0 => \N__5949\,
            in1 => \N__5906\,
            in2 => \N__5983\,
            in3 => \N__9077\,
            lcout => \uut.ir_out_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff5.q_0_neC_net\,
            ce => \N__7428\,
            sr => \_gnd_net_\
        );

    \uut.seq.q_ret_RNI52E81_0_LC_7_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__4677\,
            in1 => \N__4103\,
            in2 => \N__3803\,
            in3 => \N__4022\,
            lcout => \uut.seq.q_ret_RNI52E81Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff7.q_0_ne_LC_7_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__6388\,
            in1 => \N__6359\,
            in2 => \N__6330\,
            in3 => \N__9076\,
            lcout => \uut.ir_out_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff5.q_0_neC_net\,
            ce => \N__7428\,
            sr => \_gnd_net_\
        );

    \uut.IR.ff8.q_0_ne_LC_7_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110011111101"
        )
    port map (
            in0 => \N__9075\,
            in1 => \N__6195\,
            in2 => \N__6229\,
            in3 => \N__6885\,
            lcout => \uut.ir_out_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff5.q_0_neC_net\,
            ce => \N__7428\,
            sr => \_gnd_net_\
        );

    \uut.IR.ff3.q_RNIILCK5_LC_7_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__7987\,
            in1 => \N__7929\,
            in2 => \N__7254\,
            in3 => \N__7894\,
            lcout => OPEN,
            ltout => \uut.ir_out_m_d_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.out_1_0_iv_2_1_LC_7_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__3490\,
            in1 => \N__3436\,
            in2 => \N__3427\,
            in3 => \N__4478\,
            lcout => \uut.out_1_0_iv_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.q_ret_LC_7_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000010101010"
        )
    port map (
            in0 => \N__7406\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3884\,
            lcout => \uut.un1_HLT_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.seq.q_retC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.ALU_Out_0_7_LC_7_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001100110"
        )
    port map (
            in0 => \N__4524\,
            in1 => \N__6177\,
            in2 => \_gnd_net_\,
            in3 => \N__6768\,
            lcout => \uut.ALU_main.N_48\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.acc.ff7.q_RNIFKC71_LC_7_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6273\,
            in2 => \_gnd_net_\,
            in3 => \N__8272\,
            lcout => \uut.acc_out_m_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.out_1_0_iv_2_1_1_LC_7_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101110111"
        )
    port map (
            in0 => \N__8375\,
            in1 => \N__7247\,
            in2 => \_gnd_net_\,
            in3 => \N__7139\,
            lcout => \uut.AR_BUF.out_1_0_iv_2_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff1.q_ne_LC_7_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111110001"
        )
    port map (
            in0 => \N__9137\,
            in1 => \N__9054\,
            in2 => \N__9194\,
            in3 => \N__9239\,
            lcout => \uut.ir_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff1.q_neC_net\,
            ce => \N__7432\,
            sr => \_gnd_net_\
        );

    \uut.IR.ff2.q_ne_LC_7_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7693\,
            in1 => \N__7645\,
            in2 => \_gnd_net_\,
            in3 => \N__7597\,
            lcout => \uut.ir_out_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff1.q_neC_net\,
            ce => \N__7432\,
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_0_a5_0_2_LC_7_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__7028\,
            in1 => \N__7238\,
            in2 => \N__8716\,
            in3 => \N__4138\,
            lcout => OPEN,
            ltout => \uut.AR_BUF.g0_0_a5_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_0_a5_0_LC_7_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011000010100000"
        )
    port map (
            in0 => \N__4932\,
            in1 => \N__4702\,
            in2 => \N__3481\,
            in3 => \N__6934\,
            lcout => \uut.AR_BUF.N_9\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_1_0_1_LC_8_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110000000"
        )
    port map (
            in0 => \N__4044\,
            in1 => \N__3814\,
            in2 => \N__3469\,
            in3 => \N__3451\,
            lcout => \uut.AR_BUF.g0_1_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_0_o5_0_0_LC_8_8_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__5516\,
            in1 => \N__9402\,
            in2 => \_gnd_net_\,
            in3 => \N__8549\,
            lcout => \uut.AR_BUF.g0_0_o5_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_1_a10_3_0_LC_8_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5099\,
            in1 => \N__5357\,
            in2 => \N__3558\,
            in3 => \N__6942\,
            lcout => OPEN,
            ltout => \uut.AR_BUF.g0_1_a10_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_1_a10_LC_8_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011000000100000"
        )
    port map (
            in0 => \N__7032\,
            in1 => \N__4142\,
            in2 => \N__3454\,
            in3 => \N__4043\,
            lcout => \uut.AR_BUF.N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_1_a10_4_LC_8_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__3553\,
            in1 => \N__4930\,
            in2 => \N__3943\,
            in3 => \N__4143\,
            lcout => OPEN,
            ltout => \uut.AR_BUF.N_13_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_1_0_5_LC_8_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__5181\,
            in1 => \N__3502\,
            in2 => \N__3604\,
            in3 => \N__8253\,
            lcout => OPEN,
            ltout => \uut.AR_BUF.g0_1_0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_1_1_LC_8_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__3496\,
            in1 => \N__3565\,
            in2 => \N__3601\,
            in3 => \N__3598\,
            lcout => \uut.out_1_1_iv_3dup_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_3_a10_1_1_LC_8_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__4931\,
            in1 => \N__8757\,
            in2 => \_gnd_net_\,
            in3 => \N__5297\,
            lcout => \uut.AR_BUF.g0_3_a10_1Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_1_0_6_LC_8_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__3552\,
            in1 => \N__7760\,
            in2 => \N__3592\,
            in3 => \N__8386\,
            lcout => \uut.AR_BUF.g0_1_0_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_1_a8_3_LC_8_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__9403\,
            in1 => \N__3551\,
            in2 => \_gnd_net_\,
            in3 => \N__8550\,
            lcout => \uut.AR_BUF.N_10\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_1_0_2_LC_8_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010000000"
        )
    port map (
            in0 => \N__8577\,
            in1 => \N__8761\,
            in2 => \N__5748\,
            in3 => \N__8657\,
            lcout => \uut.AR_BUF.g0_1_0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.pc.program_counter_RNO_3_1_LC_8_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111000"
        )
    port map (
            in0 => \N__9401\,
            in1 => \N__8578\,
            in2 => \N__3664\,
            in3 => \N__7763\,
            lcout => \uut.pc.g2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.pc.program_counter_RNO_1_1_LC_8_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101011110000"
        )
    port map (
            in0 => \N__5701\,
            in1 => \_gnd_net_\,
            in2 => \N__5749\,
            in3 => \N__7327\,
            lcout => \uut.pc.N_77_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_RNICCTC1_0_LC_8_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__8656\,
            in1 => \N__5700\,
            in2 => \N__8769\,
            in3 => \N__8576\,
            lcout => \uut.program_counter_m_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.pc.program_counter_1_LC_8_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111100000"
        )
    port map (
            in0 => \N__7567\,
            in1 => \N__7643\,
            in2 => \N__5484\,
            in3 => \N__4351\,
            lcout => \uut.program_counter_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5631\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.pc.program_counter_RNO_0_0_LC_8_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000000"
        )
    port map (
            in0 => \N__9258\,
            in1 => \N__3610\,
            in2 => \N__3648\,
            in3 => \N__4207\,
            lcout => OPEN,
            ltout => \uut.pc.N_4_i_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.pc.program_counter_0_LC_8_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000011000000111"
        )
    port map (
            in0 => \N__5702\,
            in1 => \N__7328\,
            in2 => \N__3631\,
            in3 => \N__4240\,
            lcout => \uut.program_counter_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5631\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.b_reg.ff3.q_LC_8_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__8099\,
            in1 => \N__3628\,
            in2 => \N__5451\,
            in3 => \N__9053\,
            lcout => \uut.b_reg_out_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.b_reg.ff3.qC_net\,
            ce => \N__7516\,
            sr => \_gnd_net_\
        );

    \uut.ALU_main.g0_1_LC_8_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001100110"
        )
    port map (
            in0 => \N__4467\,
            in1 => \N__4499\,
            in2 => \_gnd_net_\,
            in3 => \N__6753\,
            lcout => OPEN,
            ltout => \uut.ALU_main.N_43_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_cry_1_c_RNI46ADE_LC_8_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__6581\,
            in1 => \N__6463\,
            in2 => \N__3616\,
            in3 => \N__4296\,
            lcout => \uut.alu_out_m_0_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_fast_RNIVM0N3_0_LC_8_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6752\,
            in2 => \_gnd_net_\,
            in3 => \N__4418\,
            lcout => \uut.T_1_fast_RNIVM0N3_0\,
            ltout => \uut.T_1_fast_RNIVM0N3_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.pc.program_counter_RNO_2_0_LC_8_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__6580\,
            in1 => \N__4805\,
            in2 => \N__3613\,
            in3 => \N__4320\,
            lcout => \uut.pc.N_11\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_2_rep1_RNI8TE81_LC_8_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__7020\,
            in1 => \N__4989\,
            in2 => \N__5100\,
            in3 => \N__4116\,
            lcout => OPEN,
            ltout => \uut.seq.counter.T_2_rep1_RNI8TEZ0Z81_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_2_rep1_RNI51JC1_LC_8_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3682\,
            in3 => \N__3856\,
            lcout => \uut.seq.counter.un2_MAR_LD\,
            ltout => \uut.seq.counter.un2_MAR_LD_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_RNI33MC3_3_LC_8_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__5520\,
            in1 => \N__9395\,
            in2 => \N__3679\,
            in3 => \N__8552\,
            lcout => \uut.un1_IR_OE_4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.decoder.D_0_1_LC_8_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__4990\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3855\,
            lcout => \uut.D_1_0\,
            ltout => \uut.D_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_RNIEDK31_2_LC_8_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__8744\,
            in1 => \N__4117\,
            in2 => \N__3676\,
            in3 => \N__4024\,
            lcout => \uut.un14_MAR_LD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_2_rep1_RNI6BLF1_LC_8_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111000100010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4684\,
            in2 => \_gnd_net_\,
            in3 => \N__3691\,
            lcout => \uut.T_2_rep1_RNI6BLF1\,
            ltout => \uut.T_2_rep1_RNI6BLF1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_RNIVVKI3_3_LC_8_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000100000101"
        )
    port map (
            in0 => \N__3673\,
            in1 => \N__9394\,
            in2 => \N__3667\,
            in3 => \N__8551\,
            lcout => \uut.T_1_RNIVVKI3_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.q_ret_RNI52E81_LC_8_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__4023\,
            in1 => \N__3810\,
            in2 => \N__4136\,
            in3 => \N__4685\,
            lcout => \uut.un17_IR_OE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_3_LC_8_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__8278\,
            in1 => \N__8495\,
            in2 => \N__8416\,
            in3 => \N__8359\,
            lcout => \uut.AR_BUF.g0_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff5.q_0_rep1_RNIIHI7_LC_8_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5359\,
            in2 => \_gnd_net_\,
            in3 => \N__4910\,
            lcout => OPEN,
            ltout => \uut.IR.ir_out_m_c_d_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff4.q_ne_RNINTO01_LC_8_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__8404\,
            in1 => \N__9460\,
            in2 => \N__3697\,
            in3 => \N__5082\,
            lcout => \uut.ir_out_m_c_d_3\,
            ltout => \uut.ir_out_m_c_d_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff4.q_ne_LC_8_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__9808\,
            in1 => \N__9739\,
            in2 => \N__3694\,
            in3 => \N__9859\,
            lcout => \uut.ir_out_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff4.q_neC_net\,
            ce => \N__7401\,
            sr => \_gnd_net_\
        );

    \uut.IR.ff6.q_0_ne_LC_8_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__6114\,
            in1 => \N__6141\,
            in2 => \N__9079\,
            in3 => \N__6078\,
            lcout => \uut.ir_out_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff4.q_neC_net\,
            ce => \N__7401\,
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_2_rep1_RNIGC8C1_LC_8_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__5081\,
            in1 => \N__4909\,
            in2 => \N__3733\,
            in3 => \N__4102\,
            lcout => \uut.seq.counter.T_2_rep1_RNIGC8CZ0Z1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.un13_ACC_LD_x1_LC_8_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__4982\,
            in1 => \N__4019\,
            in2 => \N__4128\,
            in3 => \N__3849\,
            lcout => OPEN,
            ltout => \uut.seq.un13_ACC_LD_xZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_fast_RNITEB42_0_LC_8_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3685\,
            in3 => \N__4839\,
            lcout => \uut.un13_ACC_LD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.decoder.D_6_LC_8_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__3731\,
            in1 => \N__5421\,
            in2 => \N__5021\,
            in3 => \N__5349\,
            lcout => \uut.D_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff7.q_ret_1_fast_LC_8_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0101010101010101"
        )
    port map (
            in0 => \N__3778\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uut.q_ret_1_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff7.q_ret_1_fastC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_2_rep1_LC_8_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7405\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uut.T_2_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff7.q_ret_1_fastC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.q_ret_RNIAFH51_LC_8_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__4020\,
            in1 => \N__3797\,
            in2 => \N__5358\,
            in3 => \N__4101\,
            lcout => \uut.un17_IR_OE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff7.q_ret_1_LC_8_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3777\,
            lcout => \uut.ir_out_i_2_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff7.q_ret_1_fastC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff7.q_0_fast_LC_8_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__4021\,
            in1 => \N__3760\,
            in2 => \_gnd_net_\,
            in3 => \N__7404\,
            lcout => \uut.q_0_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff7.q_ret_1_fastC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff5.q_0_rep1_LC_8_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7419\,
            in1 => \N__3709\,
            in2 => \_gnd_net_\,
            in3 => \N__4704\,
            lcout => \uut.ir_out_4_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff5.q_0_rep1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff8.q_0_fast_LC_8_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__3748\,
            in1 => \N__7420\,
            in2 => \_gnd_net_\,
            in3 => \N__4135\,
            lcout => \uut.q_0_fast_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff5.q_0_rep1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.decoder.D_2_0_x_LC_8_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100000000"
        )
    port map (
            in0 => \N__4978\,
            in1 => \N__5419\,
            in2 => \_gnd_net_\,
            in3 => \N__4869\,
            lcout => OPEN,
            ltout => \uut.seq.D_2_0_x_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_fast_RNI874E2_0_LC_8_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110000000000"
        )
    port map (
            in0 => \N__5012\,
            in1 => \N__4782\,
            in2 => \N__3736\,
            in3 => \N__4841\,
            lcout => \uut.S0_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff6.q_ret_1_fast_LC_8_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0011001100110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3891\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uut.q_ret_1_fast_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff5.q_0_rep1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.decoder.D_4_0_LC_8_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__5420\,
            in1 => \N__4977\,
            in2 => \N__3732\,
            in3 => \N__3848\,
            lcout => \uut.seq.D_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff5.q_0_fast_LC_8_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__7418\,
            in1 => \N__3708\,
            in2 => \_gnd_net_\,
            in3 => \N__4703\,
            lcout => \uut.ir_out_fast_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff5.q_0_rep1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_2_LC_8_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7421\,
            lcout => \uut.T_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff5.q_0_rep1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_fast_3_LC_8_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8715\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uut.seq.counter.T_1_fastZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.seq.counter.T_1_fast_3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_fast_RNI4JTR1_0_LC_8_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__7029\,
            in1 => \N__6935\,
            in2 => \N__7059\,
            in3 => \N__4843\,
            lcout => OPEN,
            ltout => \uut.seq.counter.un4_ACC_LD_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_RNI4F1C2_3_LC_8_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__9469\,
            in1 => \N__3979\,
            in2 => \N__3910\,
            in3 => \N__9396\,
            lcout => \uut.seq.counter.ACC_LD_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff6.q_ret_1_LC_8_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3892\,
            lcout => \uut.ir_out_i_2_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.seq.counter.T_1_fast_3C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_fast_RNI6J9S_3_LC_8_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011110111"
        )
    port map (
            in0 => \N__4641\,
            in1 => \N__3847\,
            in2 => \N__4988\,
            in3 => \N__9419\,
            lcout => \uut.seq.counter.T_1_fast_RNI6J9SZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_3_3_LC_9_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__4201\,
            in1 => \N__3958\,
            in2 => \N__5245\,
            in3 => \N__8286\,
            lcout => \uut.AR_BUF.g0_3Z0Z_3\,
            ltout => \uut.AR_BUF.g0_3Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.acc.ff1.q_LC_9_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011111011"
        )
    port map (
            in0 => \N__9220\,
            in1 => \N__9139\,
            in2 => \N__3826\,
            in3 => \N__9078\,
            lcout => \uut.acc_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.acc.ff1.qC_net\,
            ce => \N__5841\,
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.out_1_2_iv_1_LC_9_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__3949\,
            in1 => \N__5237\,
            in2 => \_gnd_net_\,
            in3 => \N__4200\,
            lcout => \uut.AR_BUF.out_1_2_ivZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_3_a10_0_2_LC_9_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5300\,
            in1 => \N__4144\,
            in2 => \N__8773\,
            in3 => \N__4045\,
            lcout => OPEN,
            ltout => \uut.AR_BUF.g0_3_a10_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_3_0_LC_9_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__3985\,
            in1 => \N__3978\,
            in2 => \N__3961\,
            in3 => \N__9468\,
            lcout => \uut.AR_BUF.g0_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff1.q_ne_RNIKEQ11_LC_9_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5301\,
            in2 => \_gnd_net_\,
            in3 => \N__7140\,
            lcout => OPEN,
            ltout => \uut.ir_out_m_c_d_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.out_1_2_iv_2_LC_9_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__3925\,
            in1 => \N__4225\,
            in2 => \N__3952\,
            in3 => \N__7761\,
            lcout => \uut.AR_BUF.out_1_2_ivZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_1_a10_4_1_LC_9_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5101\,
            in2 => \_gnd_net_\,
            in3 => \N__7033\,
            lcout => \uut.AR_BUF.g0_1_a10_4Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_3_2_LC_9_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110001000"
        )
    port map (
            in0 => \N__7759\,
            in1 => \N__3924\,
            in2 => \_gnd_net_\,
            in3 => \N__4224\,
            lcout => OPEN,
            ltout => \uut.AR_BUF.g0_3Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_3_6_LC_9_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111110"
        )
    port map (
            in0 => \N__5299\,
            in1 => \N__4183\,
            in2 => \N__3931\,
            in3 => \N__7893\,
            lcout => \uut.AR_BUF.g0_3Z0Z_6\,
            ltout => \uut.AR_BUF.g0_3Z0Z_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR.ff1.q_ne_LC_9_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011111011"
        )
    port map (
            in0 => \N__9175\,
            in1 => \N__9138\,
            in2 => \N__3928\,
            in3 => \N__9037\,
            lcout => \uut.AR_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.AR.ff1.q_neC_net\,
            ce => \N__8027\,
            sr => \_gnd_net_\
        );

    \uut.pc.program_counter_RNO_3_0_LC_9_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100011111111"
        )
    port map (
            in0 => \N__3923\,
            in1 => \N__7758\,
            in2 => \N__7360\,
            in3 => \N__5206\,
            lcout => OPEN,
            ltout => \uut.pc.G_26_i_a4_5_sx_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.pc.program_counter_RNO_1_0_LC_9_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__4239\,
            in1 => \N__4223\,
            in2 => \N__4210\,
            in3 => \N__4194\,
            lcout => \uut.pc.G_26_i_a4_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff1.q_ne_RNIMP2B1_LC_9_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5298\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8360\,
            lcout => \uut.ir_out_m_c_c_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_fast_RNIFJ9BG_0_LC_9_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010111000100010"
        )
    port map (
            in0 => \N__4806\,
            in1 => \N__6467\,
            in2 => \N__6603\,
            in3 => \N__4326\,
            lcout => \uut.alu_out_m_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_fast_RNIFJ9BG_0_0_LC_9_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101011001100"
        )
    port map (
            in0 => \N__4327\,
            in1 => \N__4807\,
            in2 => \N__6610\,
            in3 => \N__6474\,
            lcout => \uut.alu_out_m_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_axb_3_l_ofx_LC_9_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001101100110"
        )
    port map (
            in0 => \N__4760\,
            in1 => \N__6653\,
            in2 => \N__8497\,
            in3 => \N__4416\,
            lcout => \uut.ALU_main.un1_A_axb_3_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.b_reg.ff4.q_LC_9_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__9850\,
            in1 => \N__9802\,
            in2 => \N__9771\,
            in3 => \N__9713\,
            lcout => \uut.b_reg_out_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.b_reg.ff4.qC_net\,
            ce => \N__7487\,
            sr => \_gnd_net_\
        );

    \uut.pc.program_counter_RNO_4_1_LC_9_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001001010000000"
        )
    port map (
            in0 => \N__7549\,
            in1 => \N__6754\,
            in2 => \N__5192\,
            in3 => \N__4417\,
            lcout => OPEN,
            ltout => \uut.pc.program_counter_4_a1_0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.pc.program_counter_RNO_2_1_LC_9_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111010011110000"
        )
    port map (
            in0 => \N__6582\,
            in1 => \N__6456\,
            in2 => \N__4162\,
            in3 => \N__5124\,
            lcout => OPEN,
            ltout => \uut.pc.g1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.pc.program_counter_RNO_0_1_LC_9_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011100100"
        )
    port map (
            in0 => \N__4159\,
            in1 => \N__4153\,
            in2 => \N__4147\,
            in3 => \N__7386\,
            lcout => \uut.pc.program_counter_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_fast_RNI6RIE3_0_LC_9_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4627\,
            in2 => \_gnd_net_\,
            in3 => \N__4759\,
            lcout => \uut.un1_ALU_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_cry_0_c_THRU_CRY_0_LC_9_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4341\,
            in2 => \N__4345\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_9_12_0_\,
            carryout => \uut.ALU_main.un1_A_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_cry_0_s_LC_9_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5243\,
            in2 => \N__4534\,
            in3 => \N__4309\,
            lcout => \uut.un1_A_cry_0_s\,
            ltout => OPEN,
            carryin => \uut.ALU_main.un1_A_cry_0_c_THRU_CO\,
            carryout => \uut.ALU_main.un1_A_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_cry_0_c_RNI3CH45_LC_9_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4588\,
            in2 => \N__5193\,
            in3 => \N__4306\,
            lcout => \uut.un1_A_cry_0_c_RNI3CH45\,
            ltout => OPEN,
            carryin => \uut.ALU_main.un1_A_cry_0\,
            carryout => \uut.ALU_main.un1_A_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_cry_1_c_RNI7KL45_LC_9_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4357\,
            in2 => \N__4479\,
            in3 => \N__4285\,
            lcout => \uut.ALU_main.un1_A_cry_1_c_RNI7KLZ0Z45\,
            ltout => OPEN,
            carryin => \uut.ALU_main.un1_A_cry_1\,
            carryout => \uut.ALU_main.un1_A_cry_2_cZ0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_cry_2_c_RNIBSP45_LC_9_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4282\,
            in2 => \N__8496\,
            in3 => \N__4276\,
            lcout => \uut.un1_A_cry_2_c_RNIBSP45\,
            ltout => OPEN,
            carryin => \uut.ALU_main.un1_A_cry_2_cZ0\,
            carryout => \uut.ALU_main.un1_A_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_cry_3_c_RNIF4U45_LC_9_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4273\,
            in2 => \N__5883\,
            in3 => \N__4255\,
            lcout => \uut.ALU_main.un1_A_cry_3_c_RNIF4UZ0Z45\,
            ltout => OPEN,
            carryin => \uut.ALU_main.un1_A_cry_3\,
            carryout => \uut.ALU_main.un1_A_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_cry_4_c_RNIJC255_LC_9_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4540\,
            in2 => \N__6028\,
            in3 => \N__4243\,
            lcout => \uut.ALU_main.un1_A_cry_4_c_RNIJCZ0Z255\,
            ltout => OPEN,
            carryin => \uut.ALU_main.un1_A_cry_4\,
            carryout => \uut.ALU_main.un1_A_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_cry_5_c_RNINK655_LC_9_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4564\,
            in2 => \N__6274\,
            in3 => \N__4603\,
            lcout => \uut.ALU_main.un1_A_cry_5_c_RNINKZ0Z655\,
            ltout => OPEN,
            carryin => \uut.ALU_main.un1_A_cry_5\,
            carryout => \uut.ALU_main.un1_A_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_cry_6_c_RNINIMN4_LC_9_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4510\,
            in2 => \_gnd_net_\,
            in3 => \N__4600\,
            lcout => \uut.ALU_main.un1_A_cry_6_c_RNINIMNZ0Z4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_axb_1_l_ofx_LC_9_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100110"
        )
    port map (
            in0 => \N__7548\,
            in1 => \N__4737\,
            in2 => \N__5194\,
            in3 => \N__4396\,
            lcout => \uut.ALU_main.un1_A_axb_1_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_axb_6_l_ofx_LC_9_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010111111010"
        )
    port map (
            in0 => \N__4399\,
            in1 => \N__6265\,
            in2 => \N__4757\,
            in3 => \N__4581\,
            lcout => \uut.ALU_main.un1_A_axb_6_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_axb_5_l_ofx_LC_9_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100110"
        )
    port map (
            in0 => \N__4558\,
            in1 => \N__4739\,
            in2 => \N__6031\,
            in3 => \N__4398\,
            lcout => \uut.ALU_main.un1_A_axb_5_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_axb_0_l_ofx_LC_9_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100111100"
        )
    port map (
            in0 => \N__5244\,
            in1 => \N__6798\,
            in2 => \N__4415\,
            in3 => \N__4736\,
            lcout => \uut.ALU_main.un1_A_axb_0_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_axb_7_LC_9_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100100110110"
        )
    port map (
            in0 => \N__4400\,
            in1 => \N__4525\,
            in2 => \N__4758\,
            in3 => \N__6170\,
            lcout => \uut.ALU_main.un1_A_axbZ0Z_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_axb_2_l_ofx_LC_9_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101100110"
        )
    port map (
            in0 => \N__4504\,
            in1 => \N__4738\,
            in2 => \N__4480\,
            in3 => \N__4397\,
            lcout => \uut.ALU_main.un1_A_axb_2_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_2_rep1_RNIJDGJ_LC_9_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__5414\,
            in1 => \N__5339\,
            in2 => \N__5092\,
            in3 => \N__4906\,
            lcout => OPEN,
            ltout => \uut.seq.counter.T_2_rep1_RNIJDGJZ0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_2_rep1_RNIHU2O_LC_9_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__4786\,
            in3 => \N__4865\,
            lcout => \uut.un11_MAR_LD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.B_LD_2_tz_LC_9_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001100110011"
        )
    port map (
            in0 => \N__9458\,
            in1 => \N__4783\,
            in2 => \N__5029\,
            in3 => \N__5341\,
            lcout => \uut.B_LD_0_2_tz\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.decoder.D_0_2_LC_9_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4863\,
            in2 => \_gnd_net_\,
            in3 => \N__5413\,
            lcout => \uut.D_1_3\,
            ltout => \uut.D_1_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_fast_RNI28LI1_0_0_LC_9_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__4840\,
            in1 => \N__5340\,
            in2 => \N__4771\,
            in3 => \N__4907\,
            lcout => \uut.un7_ACC_LD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_2_rep1_RNIJ9B11_LC_9_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__5047\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5415\,
            lcout => \uut.un5_MAR_LD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.decoder.D_2_0_LC_9_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__4864\,
            in1 => \N__4981\,
            in2 => \N__5028\,
            in3 => \N__5422\,
            lcout => \uut.seq.D_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_RNIEPQK_2_LC_9_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__4908\,
            in1 => \N__4705\,
            in2 => \N__8717\,
            in3 => \N__9459\,
            lcout => \uut.un8_MAR_LD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_fast_RNIU5S31_0_LC_9_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000001"
        )
    port map (
            in0 => \N__9420\,
            in1 => \N__4642\,
            in2 => \N__5377\,
            in3 => \N__4996\,
            lcout => \uut.seq.counter.T_4\,
            ltout => \uut.seq.counter.T_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_fast_RNI4JTR1_0_0_LC_9_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111111111111"
        )
    port map (
            in0 => \N__7049\,
            in1 => \N__7019\,
            in2 => \N__4630\,
            in3 => \N__6927\,
            lcout => \uut.seq.counter.T_1_fast_RNI4JTR1_0Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_2_rep1_RNIV9NU_LC_9_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6926\,
            in1 => \N__5080\,
            in2 => \N__7031\,
            in3 => \N__4980\,
            lcout => \uut.seq.counter.T_2_rep1_RNIV9NUZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.IR.ff6.q_0_fast_LC_9_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101011001100"
        )
    port map (
            in0 => \N__5041\,
            in1 => \N__4929\,
            in2 => \_gnd_net_\,
            in3 => \N__7416\,
            lcout => \uut.q_0_fast_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff6.q_0_fastC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_fast_2_LC_9_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__7417\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uut.seq.counter.T_fastZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff6.q_0_fastC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_fast_1_LC_9_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8658\,
            lcout => \uut.seq.counter.T_1_fastZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff6.q_0_fastC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_fast_0_LC_9_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7837\,
            lcout => \uut.seq.counter.T_1_fastZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff6.q_0_fastC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.decoder.D_1_0_2_LC_9_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4979\,
            in2 => \_gnd_net_\,
            in3 => \N__5417\,
            lcout => \uut.seq.D_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.un10_ACC_LD_x1_LC_9_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__5418\,
            in1 => \N__4928\,
            in2 => \N__5356\,
            in3 => \N__4870\,
            lcout => OPEN,
            ltout => \uut.seq.un10_ACC_LD_xZ0Z1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_fast_RNI28LI1_0_LC_9_16_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110001011100010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4842\,
            in2 => \N__4813\,
            in3 => \_gnd_net_\,
            lcout => \uut.T_1_fast_RNI28LI1_0\,
            ltout => \uut.T_1_fast_RNI28LI1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.ALU_Out_0_0_LC_9_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010100001010"
        )
    port map (
            in0 => \N__5242\,
            in1 => \_gnd_net_\,
            in2 => \N__4810\,
            in3 => \N__6799\,
            lcout => \uut.N_41\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_fast_RNIH09P_2_LC_9_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__6925\,
            in1 => \N__5416\,
            in2 => \N__7030\,
            in3 => \N__5376\,
            lcout => OPEN,
            ltout => \uut.seq.counter.T_fast_RNIH09PZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_fast_RNICCPP_2_LC_9_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__5362\,
            in3 => \N__5342\,
            lcout => \uut.OUT_LD\,
            ltout => \uut.OUT_LD_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.pc.program_counter_RNO_4_0_LC_9_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100111111"
        )
    port map (
            in0 => \N__5283\,
            in1 => \N__5241\,
            in2 => \N__5209\,
            in3 => \N__7132\,
            lcout => \uut.pc.G_26_i_a4_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.ALU_Out_0_1_LC_11_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101000100"
        )
    port map (
            in0 => \N__6773\,
            in1 => \N__5182\,
            in2 => \_gnd_net_\,
            in3 => \N__7547\,
            lcout => OPEN,
            ltout => \uut.ALU_main.ALU_Out_0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_cry_0_c_RNIUP3DE_LC_11_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__6617\,
            in1 => \N__6500\,
            in2 => \N__5134\,
            in3 => \N__5131\,
            lcout => \uut.alu_out_m_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_4_LC_11_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__9393\,
            lcout => \uut.seq.counter.T_1Z0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.seq.counter.T_1_4C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.g0_0_LC_11_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001100110"
        )
    port map (
            in0 => \N__8488\,
            in1 => \N__6672\,
            in2 => \_gnd_net_\,
            in3 => \N__6772\,
            lcout => \uut.ALU_main.N_44_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_RNI215E1_0_LC_11_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5113\,
            in2 => \_gnd_net_\,
            in3 => \N__8654\,
            lcout => \uut.seq.counter.MAR_LD_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.pc.program_counter_RNO_3_3_LC_11_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__5793\,
            in1 => \N__7308\,
            in2 => \N__5763\,
            in3 => \N__5709\,
            lcout => \uut.pc.g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.pc.g0_2_LC_11_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__7309\,
            in1 => \N__5494\,
            in2 => \_gnd_net_\,
            in3 => \N__7779\,
            lcout => \uut.pc.un1_inc_0_0\,
            ltout => \uut.pc.un1_inc_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.pc.program_counter_RNO_1_3_LC_11_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5530\,
            in2 => \N__5524\,
            in3 => \N__8602\,
            lcout => \uut.pc.g0_rn_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_1_LC_11_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8655\,
            lcout => \uut.inc\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.seq.counter.T_1_1C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_RNIU1302_3_LC_11_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000100110011"
        )
    port map (
            in0 => \N__9400\,
            in1 => \N__5521\,
            in2 => \_gnd_net_\,
            in3 => \N__8574\,
            lcout => \uut.PC_LD_0_0\,
            ltout => \uut.PC_LD_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.pc.un1_inc_LC_11_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000101"
        )
    port map (
            in0 => \N__7310\,
            in1 => \_gnd_net_\,
            in2 => \N__5488\,
            in3 => \N__7780\,
            lcout => \uut.pc.un1_inc_0\,
            ltout => \uut.pc.un1_inc_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.pc.program_counter_RNO_0_2_LC_11_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000001101010011"
        )
    port map (
            in0 => \N__7209\,
            in1 => \N__5680\,
            in2 => \N__5464\,
            in3 => \N__9032\,
            lcout => \uut.pc.program_counter_4_1_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mem.data_2_7_0__m13_LC_11_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110011011"
        )
    port map (
            in0 => \N__8851\,
            in1 => \N__9607\,
            in2 => \N__9676\,
            in3 => \N__9525\,
            lcout => \uut.m13\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mar.ff2.q_ne_LC_11_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7680\,
            in1 => \N__7636\,
            in2 => \_gnd_net_\,
            in3 => \N__7589\,
            lcout => \uut.mar_out_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.mar.ff2.q_neC_net\,
            ce => \N__8799\,
            sr => \_gnd_net_\
        );

    \uut.mem.data_2_7_0__m20_LC_11_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011110111011111"
        )
    port map (
            in0 => \N__8848\,
            in1 => \N__9600\,
            in2 => \N__9675\,
            in3 => \N__9522\,
            lcout => \uut.mem.m20\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mem.data_2_7_0__m22_LC_11_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001101110111"
        )
    port map (
            in0 => \N__9524\,
            in1 => \N__9670\,
            in2 => \N__9613\,
            in3 => \N__8850\,
            lcout => \uut.mem.N_29_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mem.data_2_7_0__m18_LC_11_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011101100101"
        )
    port map (
            in0 => \N__9523\,
            in1 => \N__9671\,
            in2 => \N__9612\,
            in3 => \N__8849\,
            lcout => \uut.mem.i2_mux\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.pc.program_counter_RNO_1_2_LC_11_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101010101010"
        )
    port map (
            in0 => \N__5797\,
            in1 => \N__7311\,
            in2 => \N__5767\,
            in3 => \N__5713\,
            lcout => \uut.pc.program_counter_RNO_1Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mem.data_2_7_0__g0_0_LC_11_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110101111101111"
        )
    port map (
            in0 => \N__9520\,
            in1 => \N__8846\,
            in2 => \N__9610\,
            in3 => \N__9654\,
            lcout => \uut.N_14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.g0_LC_11_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001100110"
        )
    port map (
            in0 => \N__8464\,
            in1 => \N__6668\,
            in2 => \_gnd_net_\,
            in3 => \N__6761\,
            lcout => OPEN,
            ltout => \uut.N_44_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.pc.program_counter_RNO_0_3_LC_11_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111001001010000"
        )
    port map (
            in0 => \N__6497\,
            in1 => \N__6622\,
            in2 => \N__5674\,
            in3 => \N__6635\,
            lcout => OPEN,
            ltout => \uut.pc.alu_out_m_0_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.pc.program_counter_3_LC_11_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010101010"
        )
    port map (
            in0 => \N__5671\,
            in1 => \N__7810\,
            in2 => \N__5662\,
            in3 => \N__7843\,
            lcout => \uut.program_counter_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__5648\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mem.data_2_7_0__g0_LC_11_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010101010100000"
        )
    port map (
            in0 => \N__9521\,
            in1 => \N__8847\,
            in2 => \N__9611\,
            in3 => \N__9655\,
            lcout => \uut.N_16_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_cry_2_c_RNIAIGDE_LC_11_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__6636\,
            in1 => \N__6614\,
            in2 => \N__5542\,
            in3 => \N__6498\,
            lcout => \uut.alu_out_m_1_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.ALU_Out_0_3_LC_11_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010010101010000"
        )
    port map (
            in0 => \N__6762\,
            in1 => \_gnd_net_\,
            in2 => \N__6673\,
            in3 => \N__8465\,
            lcout => OPEN,
            ltout => \uut.ALU_main.N_44_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.ALU_main.un1_A_cry_2_c_RNIAIGDE_0_LC_11_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__6637\,
            in1 => \N__6615\,
            in2 => \N__6505\,
            in3 => \N__6499\,
            lcout => \uut.alu_out_m_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.acc.ff4.q_LC_11_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__9804\,
            in1 => \N__9852\,
            in2 => \N__9763\,
            in3 => \N__9718\,
            lcout => \uut.acc_out_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.acc.ff4.qC_net\,
            ce => \N__5837\,
            sr => \_gnd_net_\
        );

    \uut.acc.ff7.q_LC_11_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__6406\,
            in1 => \N__6367\,
            in2 => \N__6320\,
            in3 => \N__8975\,
            lcout => \uut.acc_out_6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.acc.ff4.qC_net\,
            ce => \N__5837\,
            sr => \_gnd_net_\
        );

    \uut.acc.ff8.q_LC_11_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001101"
        )
    port map (
            in0 => \N__8972\,
            in1 => \N__6228\,
            in2 => \N__6884\,
            in3 => \N__6199\,
            lcout => \uut.acc_out_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.acc.ff4.qC_net\,
            ce => \N__5837\,
            sr => \_gnd_net_\
        );

    \uut.acc.ff6.q_LC_11_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__6145\,
            in1 => \N__6115\,
            in2 => \N__6070\,
            in3 => \N__8974\,
            lcout => \uut.acc_out_5\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.acc.ff4.qC_net\,
            ce => \N__5837\,
            sr => \_gnd_net_\
        );

    \uut.acc.ff5.q_LC_11_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111001101"
        )
    port map (
            in0 => \N__8973\,
            in1 => \N__5979\,
            in2 => \N__5953\,
            in3 => \N__5917\,
            lcout => \uut.acc_out_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.acc.ff4.qC_net\,
            ce => \N__5837\,
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_RNIFRTJ2_3_LC_11_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011001100"
        )
    port map (
            in0 => \N__9279\,
            in1 => \N__9363\,
            in2 => \_gnd_net_\,
            in3 => \N__9310\,
            lcout => \uut.B_LD_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.B_LD_1_tz_LC_11_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__7060\,
            in1 => \N__7027\,
            in2 => \N__6955\,
            in3 => \N__6943\,
            lcout => \uut.B_LD_0_1_tz\,
            ltout => \uut.B_LD_0_1_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_RNII3T14_3_LC_11_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1011001100000000"
        )
    port map (
            in0 => \N__9278\,
            in1 => \N__9362\,
            in2 => \N__6892\,
            in3 => \N__9297\,
            lcout => \uut.ROM_OE\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mem.data_2_7_0__m26_LC_11_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111011001101101"
        )
    port map (
            in0 => \N__8843\,
            in1 => \N__9589\,
            in2 => \N__9544\,
            in3 => \N__9653\,
            lcout => \uut.mem.i2_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.out_reg.ff3.q_LC_11_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011110000"
        )
    port map (
            in0 => \N__8077\,
            in1 => \N__6847\,
            in2 => \N__6834\,
            in3 => \N__8280\,
            lcout => \LED3_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.out_reg.ff3.qC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_3_LC_11_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8768\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \uut.T_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.out_reg.ff3.qC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mem.data_2_7_0__m10_LC_11_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111001111"
        )
    port map (
            in0 => \N__9652\,
            in1 => \N__9539\,
            in2 => \N__9608\,
            in3 => \N__8842\,
            lcout => \uut.m10\,
            ltout => \uut.m10_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mem.data_2_7_0__N_11_i_m_LC_11_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6802\,
            in3 => \N__8923\,
            lcout => \uut.N_11_i_m\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.b_reg.ff1.q_LC_11_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011111011"
        )
    port map (
            in0 => \N__9240\,
            in1 => \N__9123\,
            in2 => \N__9195\,
            in3 => \N__8976\,
            lcout => \uut.b_reg_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.b_reg.ff1.qC_net\,
            ce => \N__7481\,
            sr => \_gnd_net_\
        );

    \uut.b_reg.ff2.q_LC_11_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111101110"
        )
    port map (
            in0 => \N__7688\,
            in1 => \N__7623\,
            in2 => \_gnd_net_\,
            in3 => \N__7596\,
            lcout => \uut.b_reg_out_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.b_reg.ff1.qC_net\,
            ce => \N__7481\,
            sr => \_gnd_net_\
        );

    \uut.IR.ff3.q_LC_11_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111101011001100"
        )
    port map (
            in0 => \N__8073\,
            in1 => \N__7237\,
            in2 => \N__8125\,
            in3 => \N__7402\,
            lcout => \uut.ir_out_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.IR.ff3.qC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_RNI3K4S_2_LC_12_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__8575\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8767\,
            lcout => \uut.AR_LD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_9_LC_12_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111100010001"
        )
    port map (
            in0 => \N__7210\,
            in1 => \N__9033\,
            in2 => \_gnd_net_\,
            in3 => \N__7192\,
            lcout => \uut.out_1_0_iv_3\,
            ltout => \uut.out_1_0_iv_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR.ff3.q_LC_12_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110110101000"
        )
    port map (
            in0 => \N__8023\,
            in1 => \N__8108\,
            in2 => \N__7174\,
            in3 => \N__7163\,
            lcout => \uut.AR_out_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.AR.ff3.qC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_2_rep1_RNI48EP1_LC_12_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8384\,
            in2 => \_gnd_net_\,
            in3 => \N__7141\,
            lcout => \uut.MAR_LD_1\,
            ltout => \uut.MAR_LD_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_RNI2G205_0_LC_12_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100000"
        )
    port map (
            in0 => \N__7090\,
            in1 => \N__7986\,
            in2 => \N__7084\,
            in3 => \N__7939\,
            lcout => \uut.MAR_LD_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_5_LC_12_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001101"
        )
    port map (
            in0 => \N__8985\,
            in1 => \N__7699\,
            in2 => \N__7081\,
            in3 => \N__7072\,
            lcout => \uut.AR_BUF.g0Z0Z_5\,
            ltout => \uut.AR_BUF.g0Z0Z_5_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR.ff4.q_ne_LC_12_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__9712\,
            in1 => \N__9767\,
            in2 => \N__7063\,
            in3 => \N__9836\,
            lcout => \uut.AR_out_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.AR.ff4.q_neC_net\,
            ce => \N__8031\,
            sr => \_gnd_net_\
        );

    \uut.IR.ff4.q_ne_RNI59RD5_LC_12_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011110000"
        )
    port map (
            in0 => \N__7985\,
            in1 => \N__7935\,
            in2 => \N__8431\,
            in3 => \N__7892\,
            lcout => \uut.ir_out_m_d_3\,
            ltout => \uut.ir_out_m_d_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.pc.program_counter_RNO_2_3_LC_12_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__7852\,
            in2 => \N__7846\,
            in3 => \N__8301\,
            lcout => \uut.pc.g0_sn\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.out_1_iv_2_LC_12_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__8503\,
            in1 => \N__9711\,
            in2 => \N__7803\,
            in3 => \N__7781\,
            lcout => \uut.out_1_iv_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_0_LC_12_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7836\,
            lcout => \uut.T_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.seq.counter.T_1_0C_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.out_1_ivdup_0_LC_12_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__8261\,
            in1 => \N__8426\,
            in2 => \N__8478\,
            in3 => \N__8383\,
            lcout => OPEN,
            ltout => \uut.AR_BUF.out_1_ivdupZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_0_LC_12_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000011110111"
        )
    port map (
            in0 => \N__9865\,
            in1 => \N__9526\,
            in2 => \N__7813\,
            in3 => \N__8984\,
            lcout => \uut.g0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_RNI0KMT_0_LC_12_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011001100"
        )
    port map (
            in0 => \N__8766\,
            in1 => \N__8634\,
            in2 => \_gnd_net_\,
            in3 => \N__8581\,
            lcout => OPEN,
            ltout => \uut.g1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.g0_2_LC_12_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__7804\,
            in1 => \N__8597\,
            in2 => \N__7786\,
            in3 => \N__7782\,
            lcout => \uut.AR_BUF.g0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_RNIFFTC1_0_LC_12_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110000011000000"
        )
    port map (
            in0 => \N__8765\,
            in1 => \N__8633\,
            in2 => \N__8601\,
            in3 => \N__8580\,
            lcout => \uut.program_counter_m_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.out_1_iv_0_LC_12_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111010101010"
        )
    port map (
            in0 => \N__8477\,
            in1 => \N__8430\,
            in2 => \_gnd_net_\,
            in3 => \N__8382\,
            lcout => OPEN,
            ltout => \uut.AR_BUF.out_1_ivZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.out_1_iv_2_1_LC_12_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__9840\,
            in2 => \N__8308\,
            in3 => \N__8305\,
            lcout => OPEN,
            ltout => \uut.out_1_iv_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.out_reg.ff4.q_LC_12_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111110010101010"
        )
    port map (
            in0 => \N__8157\,
            in1 => \N__8131\,
            in2 => \N__8290\,
            in3 => \N__8279\,
            lcout => \LED4_c\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.out_reg.ff4.qC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mem.data_2_7_0__m15_LC_12_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100011001000"
        )
    port map (
            in0 => \N__9665\,
            in1 => \N__9535\,
            in2 => \N__9609\,
            in3 => \N__8845\,
            lcout => OPEN,
            ltout => \uut.m15_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.AR_BUF.out_1_iv_3_LC_12_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8140\,
            in2 => \N__8134\,
            in3 => \N__8971\,
            lcout => \uut.out_1_iv_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mar.ff1.q_sbtinv_LC_12_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8043\,
            lcout => \uut.mar.MAR_LD_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mar.ff3.q_LC_12_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111000001110"
        )
    port map (
            in0 => \N__8121\,
            in1 => \N__8066\,
            in2 => \N__8047\,
            in3 => \N__9666\,
            lcout => \uut.mar_out_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.out_reg.ff4.qC_net\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mem.data_2_7_0__g1_LC_12_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011101110"
        )
    port map (
            in0 => \N__9590\,
            in1 => \N__9651\,
            in2 => \_gnd_net_\,
            in3 => \N__8844\,
            lcout => \uut.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mar.ff4.q_ne_LC_12_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1111111111111110"
        )
    port map (
            in0 => \N__9851\,
            in1 => \N__9803\,
            in2 => \N__9772\,
            in3 => \N__9714\,
            lcout => \uut.mar_out_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.mar.ff4.q_neC_net\,
            ce => \N__8800\,
            sr => \_gnd_net_\
        );

    \uut.mem.data_2_7_0__m6_LC_12_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110100111"
        )
    port map (
            in0 => \N__9650\,
            in1 => \N__9571\,
            in2 => \N__9543\,
            in3 => \N__8827\,
            lcout => \uut.m6\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.seq.counter.T_1_fast_RNI38VD1_1_LC_12_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010111011"
        )
    port map (
            in0 => \N__9481\,
            in1 => \N__9464\,
            in2 => \_gnd_net_\,
            in3 => \N__9427\,
            lcout => \uut.un1_ROM_OE_0\,
            ltout => \uut.un1_ROM_OE_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mem.data_2_7_0__N_7_i_m_sx_LC_12_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101010000"
        )
    port map (
            in0 => \N__9356\,
            in1 => \_gnd_net_\,
            in2 => \N__9313\,
            in3 => \N__9110\,
            lcout => OPEN,
            ltout => \uut.mem.N_7_i_m_sx_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mem.data_2_7_0__N_7_i_m_LC_12_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__9309\,
            in1 => \N__9298\,
            in2 => \N__9286\,
            in3 => \N__9283\,
            lcout => \uut.N_7_i_m\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \uut.mar.ff1.q_ne_LC_12_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__9241\,
            in1 => \N__9196\,
            in2 => \N__9133\,
            in3 => \N__8977\,
            lcout => \uut.mar_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVuut.mar.ff4.q_neC_net\,
            ce => \N__8800\,
            sr => \_gnd_net_\
        );
end \INTERFACE\;
