// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Dec 13 2023 18:09:27

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "main" view "INTERFACE"

module main (
    out,
    clr,
    clk);

    output [7:0] out;
    input clr;
    input clk;

    wire N__9029;
    wire N__9028;
    wire N__9027;
    wire N__9018;
    wire N__9017;
    wire N__9016;
    wire N__9009;
    wire N__9008;
    wire N__9007;
    wire N__9000;
    wire N__8999;
    wire N__8998;
    wire N__8991;
    wire N__8990;
    wire N__8989;
    wire N__8982;
    wire N__8981;
    wire N__8980;
    wire N__8973;
    wire N__8972;
    wire N__8971;
    wire N__8964;
    wire N__8963;
    wire N__8962;
    wire N__8955;
    wire N__8954;
    wire N__8953;
    wire N__8946;
    wire N__8945;
    wire N__8944;
    wire N__8927;
    wire N__8926;
    wire N__8923;
    wire N__8920;
    wire N__8919;
    wire N__8916;
    wire N__8913;
    wire N__8910;
    wire N__8909;
    wire N__8908;
    wire N__8901;
    wire N__8898;
    wire N__8895;
    wire N__8892;
    wire N__8889;
    wire N__8886;
    wire N__8879;
    wire N__8878;
    wire N__8877;
    wire N__8874;
    wire N__8873;
    wire N__8870;
    wire N__8867;
    wire N__8864;
    wire N__8861;
    wire N__8860;
    wire N__8857;
    wire N__8854;
    wire N__8849;
    wire N__8848;
    wire N__8845;
    wire N__8842;
    wire N__8839;
    wire N__8836;
    wire N__8833;
    wire N__8830;
    wire N__8825;
    wire N__8816;
    wire N__8815;
    wire N__8814;
    wire N__8811;
    wire N__8808;
    wire N__8807;
    wire N__8804;
    wire N__8799;
    wire N__8796;
    wire N__8795;
    wire N__8794;
    wire N__8791;
    wire N__8788;
    wire N__8785;
    wire N__8782;
    wire N__8779;
    wire N__8776;
    wire N__8765;
    wire N__8764;
    wire N__8763;
    wire N__8760;
    wire N__8757;
    wire N__8756;
    wire N__8755;
    wire N__8752;
    wire N__8749;
    wire N__8748;
    wire N__8745;
    wire N__8742;
    wire N__8739;
    wire N__8736;
    wire N__8733;
    wire N__8732;
    wire N__8731;
    wire N__8728;
    wire N__8723;
    wire N__8720;
    wire N__8715;
    wire N__8712;
    wire N__8709;
    wire N__8706;
    wire N__8703;
    wire N__8698;
    wire N__8687;
    wire N__8686;
    wire N__8685;
    wire N__8684;
    wire N__8683;
    wire N__8680;
    wire N__8679;
    wire N__8678;
    wire N__8677;
    wire N__8676;
    wire N__8675;
    wire N__8674;
    wire N__8673;
    wire N__8672;
    wire N__8669;
    wire N__8668;
    wire N__8667;
    wire N__8666;
    wire N__8665;
    wire N__8664;
    wire N__8663;
    wire N__8662;
    wire N__8661;
    wire N__8660;
    wire N__8659;
    wire N__8656;
    wire N__8655;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8645;
    wire N__8642;
    wire N__8639;
    wire N__8636;
    wire N__8633;
    wire N__8630;
    wire N__8625;
    wire N__8622;
    wire N__8621;
    wire N__8614;
    wire N__8609;
    wire N__8604;
    wire N__8601;
    wire N__8596;
    wire N__8587;
    wire N__8584;
    wire N__8579;
    wire N__8576;
    wire N__8573;
    wire N__8568;
    wire N__8563;
    wire N__8560;
    wire N__8557;
    wire N__8554;
    wire N__8553;
    wire N__8552;
    wire N__8551;
    wire N__8550;
    wire N__8549;
    wire N__8548;
    wire N__8545;
    wire N__8534;
    wire N__8531;
    wire N__8528;
    wire N__8523;
    wire N__8514;
    wire N__8509;
    wire N__8500;
    wire N__8495;
    wire N__8480;
    wire N__8479;
    wire N__8478;
    wire N__8475;
    wire N__8472;
    wire N__8469;
    wire N__8468;
    wire N__8461;
    wire N__8458;
    wire N__8457;
    wire N__8452;
    wire N__8449;
    wire N__8448;
    wire N__8443;
    wire N__8440;
    wire N__8435;
    wire N__8434;
    wire N__8431;
    wire N__8428;
    wire N__8427;
    wire N__8426;
    wire N__8425;
    wire N__8422;
    wire N__8419;
    wire N__8416;
    wire N__8413;
    wire N__8412;
    wire N__8411;
    wire N__8408;
    wire N__8403;
    wire N__8400;
    wire N__8397;
    wire N__8394;
    wire N__8391;
    wire N__8386;
    wire N__8375;
    wire N__8374;
    wire N__8373;
    wire N__8370;
    wire N__8369;
    wire N__8368;
    wire N__8365;
    wire N__8362;
    wire N__8359;
    wire N__8356;
    wire N__8353;
    wire N__8350;
    wire N__8347;
    wire N__8344;
    wire N__8341;
    wire N__8338;
    wire N__8335;
    wire N__8332;
    wire N__8325;
    wire N__8322;
    wire N__8319;
    wire N__8316;
    wire N__8309;
    wire N__8308;
    wire N__8307;
    wire N__8306;
    wire N__8303;
    wire N__8300;
    wire N__8297;
    wire N__8294;
    wire N__8293;
    wire N__8290;
    wire N__8283;
    wire N__8280;
    wire N__8279;
    wire N__8272;
    wire N__8269;
    wire N__8266;
    wire N__8263;
    wire N__8258;
    wire N__8257;
    wire N__8254;
    wire N__8253;
    wire N__8246;
    wire N__8243;
    wire N__8240;
    wire N__8237;
    wire N__8236;
    wire N__8233;
    wire N__8230;
    wire N__8229;
    wire N__8228;
    wire N__8223;
    wire N__8220;
    wire N__8217;
    wire N__8212;
    wire N__8211;
    wire N__8210;
    wire N__8207;
    wire N__8204;
    wire N__8201;
    wire N__8198;
    wire N__8193;
    wire N__8188;
    wire N__8183;
    wire N__8182;
    wire N__8179;
    wire N__8176;
    wire N__8173;
    wire N__8170;
    wire N__8169;
    wire N__8168;
    wire N__8167;
    wire N__8166;
    wire N__8161;
    wire N__8158;
    wire N__8155;
    wire N__8152;
    wire N__8149;
    wire N__8138;
    wire N__8137;
    wire N__8134;
    wire N__8131;
    wire N__8130;
    wire N__8129;
    wire N__8126;
    wire N__8123;
    wire N__8122;
    wire N__8121;
    wire N__8118;
    wire N__8115;
    wire N__8114;
    wire N__8109;
    wire N__8106;
    wire N__8103;
    wire N__8100;
    wire N__8097;
    wire N__8094;
    wire N__8091;
    wire N__8088;
    wire N__8085;
    wire N__8080;
    wire N__8077;
    wire N__8066;
    wire N__8065;
    wire N__8064;
    wire N__8061;
    wire N__8060;
    wire N__8057;
    wire N__8054;
    wire N__8053;
    wire N__8052;
    wire N__8049;
    wire N__8046;
    wire N__8045;
    wire N__8042;
    wire N__8039;
    wire N__8036;
    wire N__8033;
    wire N__8028;
    wire N__8025;
    wire N__8012;
    wire N__8009;
    wire N__8006;
    wire N__8003;
    wire N__8002;
    wire N__7999;
    wire N__7996;
    wire N__7995;
    wire N__7994;
    wire N__7991;
    wire N__7988;
    wire N__7985;
    wire N__7982;
    wire N__7977;
    wire N__7974;
    wire N__7971;
    wire N__7964;
    wire N__7961;
    wire N__7960;
    wire N__7959;
    wire N__7956;
    wire N__7953;
    wire N__7952;
    wire N__7951;
    wire N__7948;
    wire N__7945;
    wire N__7942;
    wire N__7939;
    wire N__7936;
    wire N__7933;
    wire N__7922;
    wire N__7919;
    wire N__7916;
    wire N__7915;
    wire N__7914;
    wire N__7911;
    wire N__7910;
    wire N__7909;
    wire N__7908;
    wire N__7905;
    wire N__7904;
    wire N__7903;
    wire N__7900;
    wire N__7897;
    wire N__7892;
    wire N__7889;
    wire N__7886;
    wire N__7883;
    wire N__7878;
    wire N__7873;
    wire N__7870;
    wire N__7867;
    wire N__7864;
    wire N__7857;
    wire N__7854;
    wire N__7849;
    wire N__7844;
    wire N__7841;
    wire N__7838;
    wire N__7835;
    wire N__7834;
    wire N__7833;
    wire N__7830;
    wire N__7825;
    wire N__7822;
    wire N__7819;
    wire N__7816;
    wire N__7811;
    wire N__7808;
    wire N__7805;
    wire N__7804;
    wire N__7803;
    wire N__7800;
    wire N__7797;
    wire N__7794;
    wire N__7793;
    wire N__7788;
    wire N__7785;
    wire N__7782;
    wire N__7781;
    wire N__7778;
    wire N__7773;
    wire N__7770;
    wire N__7767;
    wire N__7764;
    wire N__7761;
    wire N__7754;
    wire N__7751;
    wire N__7750;
    wire N__7749;
    wire N__7748;
    wire N__7745;
    wire N__7742;
    wire N__7741;
    wire N__7740;
    wire N__7737;
    wire N__7734;
    wire N__7729;
    wire N__7726;
    wire N__7723;
    wire N__7720;
    wire N__7717;
    wire N__7714;
    wire N__7711;
    wire N__7706;
    wire N__7703;
    wire N__7700;
    wire N__7697;
    wire N__7694;
    wire N__7685;
    wire N__7682;
    wire N__7681;
    wire N__7680;
    wire N__7679;
    wire N__7678;
    wire N__7675;
    wire N__7672;
    wire N__7669;
    wire N__7666;
    wire N__7663;
    wire N__7660;
    wire N__7657;
    wire N__7654;
    wire N__7649;
    wire N__7646;
    wire N__7643;
    wire N__7638;
    wire N__7631;
    wire N__7630;
    wire N__7627;
    wire N__7624;
    wire N__7621;
    wire N__7620;
    wire N__7619;
    wire N__7618;
    wire N__7615;
    wire N__7612;
    wire N__7609;
    wire N__7606;
    wire N__7603;
    wire N__7600;
    wire N__7597;
    wire N__7594;
    wire N__7593;
    wire N__7590;
    wire N__7587;
    wire N__7584;
    wire N__7579;
    wire N__7576;
    wire N__7573;
    wire N__7570;
    wire N__7567;
    wire N__7564;
    wire N__7561;
    wire N__7556;
    wire N__7547;
    wire N__7546;
    wire N__7545;
    wire N__7544;
    wire N__7541;
    wire N__7540;
    wire N__7537;
    wire N__7534;
    wire N__7531;
    wire N__7528;
    wire N__7525;
    wire N__7524;
    wire N__7521;
    wire N__7518;
    wire N__7515;
    wire N__7510;
    wire N__7507;
    wire N__7500;
    wire N__7493;
    wire N__7490;
    wire N__7487;
    wire N__7484;
    wire N__7481;
    wire N__7480;
    wire N__7479;
    wire N__7478;
    wire N__7477;
    wire N__7476;
    wire N__7475;
    wire N__7474;
    wire N__7473;
    wire N__7470;
    wire N__7467;
    wire N__7464;
    wire N__7461;
    wire N__7458;
    wire N__7457;
    wire N__7456;
    wire N__7455;
    wire N__7454;
    wire N__7451;
    wire N__7448;
    wire N__7445;
    wire N__7442;
    wire N__7441;
    wire N__7438;
    wire N__7435;
    wire N__7432;
    wire N__7427;
    wire N__7424;
    wire N__7419;
    wire N__7416;
    wire N__7413;
    wire N__7412;
    wire N__7409;
    wire N__7404;
    wire N__7401;
    wire N__7400;
    wire N__7399;
    wire N__7398;
    wire N__7389;
    wire N__7388;
    wire N__7385;
    wire N__7378;
    wire N__7375;
    wire N__7370;
    wire N__7367;
    wire N__7364;
    wire N__7361;
    wire N__7358;
    wire N__7355;
    wire N__7352;
    wire N__7345;
    wire N__7340;
    wire N__7333;
    wire N__7322;
    wire N__7321;
    wire N__7320;
    wire N__7319;
    wire N__7318;
    wire N__7317;
    wire N__7316;
    wire N__7315;
    wire N__7314;
    wire N__7313;
    wire N__7312;
    wire N__7311;
    wire N__7310;
    wire N__7309;
    wire N__7308;
    wire N__7307;
    wire N__7306;
    wire N__7305;
    wire N__7304;
    wire N__7303;
    wire N__7302;
    wire N__7301;
    wire N__7300;
    wire N__7299;
    wire N__7298;
    wire N__7297;
    wire N__7296;
    wire N__7295;
    wire N__7294;
    wire N__7293;
    wire N__7292;
    wire N__7291;
    wire N__7290;
    wire N__7289;
    wire N__7288;
    wire N__7287;
    wire N__7214;
    wire N__7211;
    wire N__7208;
    wire N__7205;
    wire N__7202;
    wire N__7199;
    wire N__7196;
    wire N__7193;
    wire N__7192;
    wire N__7187;
    wire N__7186;
    wire N__7183;
    wire N__7180;
    wire N__7179;
    wire N__7178;
    wire N__7177;
    wire N__7176;
    wire N__7175;
    wire N__7174;
    wire N__7173;
    wire N__7168;
    wire N__7167;
    wire N__7156;
    wire N__7151;
    wire N__7148;
    wire N__7145;
    wire N__7142;
    wire N__7139;
    wire N__7130;
    wire N__7129;
    wire N__7128;
    wire N__7127;
    wire N__7122;
    wire N__7121;
    wire N__7120;
    wire N__7119;
    wire N__7118;
    wire N__7115;
    wire N__7114;
    wire N__7113;
    wire N__7110;
    wire N__7109;
    wire N__7108;
    wire N__7105;
    wire N__7102;
    wire N__7099;
    wire N__7094;
    wire N__7083;
    wire N__7080;
    wire N__7077;
    wire N__7070;
    wire N__7067;
    wire N__7058;
    wire N__7057;
    wire N__7054;
    wire N__7053;
    wire N__7048;
    wire N__7047;
    wire N__7046;
    wire N__7045;
    wire N__7044;
    wire N__7043;
    wire N__7042;
    wire N__7039;
    wire N__7036;
    wire N__7033;
    wire N__7030;
    wire N__7029;
    wire N__7028;
    wire N__7025;
    wire N__7022;
    wire N__7019;
    wire N__7018;
    wire N__7015;
    wire N__7012;
    wire N__7009;
    wire N__6998;
    wire N__6995;
    wire N__6988;
    wire N__6985;
    wire N__6980;
    wire N__6975;
    wire N__6968;
    wire N__6967;
    wire N__6966;
    wire N__6965;
    wire N__6964;
    wire N__6963;
    wire N__6962;
    wire N__6961;
    wire N__6960;
    wire N__6957;
    wire N__6952;
    wire N__6949;
    wire N__6938;
    wire N__6935;
    wire N__6934;
    wire N__6933;
    wire N__6932;
    wire N__6927;
    wire N__6924;
    wire N__6921;
    wire N__6914;
    wire N__6909;
    wire N__6902;
    wire N__6901;
    wire N__6900;
    wire N__6895;
    wire N__6892;
    wire N__6891;
    wire N__6890;
    wire N__6887;
    wire N__6884;
    wire N__6881;
    wire N__6878;
    wire N__6875;
    wire N__6872;
    wire N__6869;
    wire N__6866;
    wire N__6863;
    wire N__6854;
    wire N__6851;
    wire N__6848;
    wire N__6847;
    wire N__6844;
    wire N__6841;
    wire N__6836;
    wire N__6833;
    wire N__6830;
    wire N__6829;
    wire N__6826;
    wire N__6823;
    wire N__6822;
    wire N__6821;
    wire N__6820;
    wire N__6817;
    wire N__6814;
    wire N__6811;
    wire N__6808;
    wire N__6805;
    wire N__6800;
    wire N__6791;
    wire N__6790;
    wire N__6789;
    wire N__6786;
    wire N__6783;
    wire N__6782;
    wire N__6779;
    wire N__6778;
    wire N__6775;
    wire N__6772;
    wire N__6769;
    wire N__6766;
    wire N__6763;
    wire N__6756;
    wire N__6753;
    wire N__6746;
    wire N__6745;
    wire N__6742;
    wire N__6739;
    wire N__6736;
    wire N__6735;
    wire N__6734;
    wire N__6729;
    wire N__6726;
    wire N__6723;
    wire N__6720;
    wire N__6717;
    wire N__6714;
    wire N__6711;
    wire N__6704;
    wire N__6703;
    wire N__6700;
    wire N__6697;
    wire N__6692;
    wire N__6691;
    wire N__6690;
    wire N__6687;
    wire N__6684;
    wire N__6683;
    wire N__6680;
    wire N__6677;
    wire N__6674;
    wire N__6671;
    wire N__6670;
    wire N__6667;
    wire N__6664;
    wire N__6661;
    wire N__6658;
    wire N__6655;
    wire N__6652;
    wire N__6641;
    wire N__6638;
    wire N__6637;
    wire N__6636;
    wire N__6635;
    wire N__6634;
    wire N__6631;
    wire N__6628;
    wire N__6625;
    wire N__6622;
    wire N__6619;
    wire N__6610;
    wire N__6605;
    wire N__6604;
    wire N__6601;
    wire N__6600;
    wire N__6599;
    wire N__6598;
    wire N__6595;
    wire N__6592;
    wire N__6589;
    wire N__6586;
    wire N__6583;
    wire N__6580;
    wire N__6575;
    wire N__6572;
    wire N__6569;
    wire N__6564;
    wire N__6557;
    wire N__6556;
    wire N__6555;
    wire N__6554;
    wire N__6553;
    wire N__6552;
    wire N__6551;
    wire N__6548;
    wire N__6543;
    wire N__6538;
    wire N__6537;
    wire N__6536;
    wire N__6535;
    wire N__6534;
    wire N__6531;
    wire N__6528;
    wire N__6527;
    wire N__6526;
    wire N__6525;
    wire N__6524;
    wire N__6523;
    wire N__6522;
    wire N__6521;
    wire N__6514;
    wire N__6511;
    wire N__6504;
    wire N__6499;
    wire N__6496;
    wire N__6489;
    wire N__6486;
    wire N__6483;
    wire N__6482;
    wire N__6479;
    wire N__6474;
    wire N__6467;
    wire N__6466;
    wire N__6465;
    wire N__6464;
    wire N__6463;
    wire N__6460;
    wire N__6455;
    wire N__6452;
    wire N__6445;
    wire N__6438;
    wire N__6435;
    wire N__6422;
    wire N__6419;
    wire N__6416;
    wire N__6413;
    wire N__6410;
    wire N__6407;
    wire N__6404;
    wire N__6401;
    wire N__6398;
    wire N__6395;
    wire N__6392;
    wire N__6389;
    wire N__6386;
    wire N__6383;
    wire N__6382;
    wire N__6379;
    wire N__6376;
    wire N__6373;
    wire N__6370;
    wire N__6365;
    wire N__6362;
    wire N__6359;
    wire N__6358;
    wire N__6353;
    wire N__6350;
    wire N__6347;
    wire N__6346;
    wire N__6343;
    wire N__6340;
    wire N__6335;
    wire N__6334;
    wire N__6331;
    wire N__6328;
    wire N__6327;
    wire N__6324;
    wire N__6321;
    wire N__6318;
    wire N__6311;
    wire N__6310;
    wire N__6309;
    wire N__6306;
    wire N__6303;
    wire N__6300;
    wire N__6297;
    wire N__6294;
    wire N__6293;
    wire N__6290;
    wire N__6285;
    wire N__6282;
    wire N__6279;
    wire N__6276;
    wire N__6269;
    wire N__6268;
    wire N__6265;
    wire N__6262;
    wire N__6259;
    wire N__6256;
    wire N__6251;
    wire N__6248;
    wire N__6245;
    wire N__6244;
    wire N__6243;
    wire N__6240;
    wire N__6235;
    wire N__6232;
    wire N__6229;
    wire N__6224;
    wire N__6221;
    wire N__6218;
    wire N__6215;
    wire N__6212;
    wire N__6209;
    wire N__6206;
    wire N__6205;
    wire N__6202;
    wire N__6199;
    wire N__6194;
    wire N__6193;
    wire N__6192;
    wire N__6191;
    wire N__6190;
    wire N__6187;
    wire N__6186;
    wire N__6183;
    wire N__6180;
    wire N__6175;
    wire N__6172;
    wire N__6169;
    wire N__6168;
    wire N__6167;
    wire N__6166;
    wire N__6165;
    wire N__6164;
    wire N__6163;
    wire N__6162;
    wire N__6161;
    wire N__6160;
    wire N__6159;
    wire N__6158;
    wire N__6157;
    wire N__6156;
    wire N__6153;
    wire N__6148;
    wire N__6143;
    wire N__6136;
    wire N__6131;
    wire N__6124;
    wire N__6119;
    wire N__6112;
    wire N__6095;
    wire N__6092;
    wire N__6089;
    wire N__6086;
    wire N__6083;
    wire N__6080;
    wire N__6079;
    wire N__6076;
    wire N__6073;
    wire N__6068;
    wire N__6067;
    wire N__6064;
    wire N__6061;
    wire N__6060;
    wire N__6055;
    wire N__6052;
    wire N__6051;
    wire N__6050;
    wire N__6045;
    wire N__6042;
    wire N__6039;
    wire N__6036;
    wire N__6029;
    wire N__6028;
    wire N__6025;
    wire N__6024;
    wire N__6021;
    wire N__6018;
    wire N__6015;
    wire N__6014;
    wire N__6011;
    wire N__6006;
    wire N__6003;
    wire N__6000;
    wire N__5993;
    wire N__5992;
    wire N__5991;
    wire N__5990;
    wire N__5989;
    wire N__5986;
    wire N__5979;
    wire N__5976;
    wire N__5973;
    wire N__5970;
    wire N__5967;
    wire N__5964;
    wire N__5961;
    wire N__5958;
    wire N__5955;
    wire N__5948;
    wire N__5947;
    wire N__5944;
    wire N__5941;
    wire N__5938;
    wire N__5935;
    wire N__5932;
    wire N__5929;
    wire N__5924;
    wire N__5921;
    wire N__5918;
    wire N__5915;
    wire N__5912;
    wire N__5909;
    wire N__5908;
    wire N__5907;
    wire N__5906;
    wire N__5903;
    wire N__5900;
    wire N__5895;
    wire N__5892;
    wire N__5885;
    wire N__5882;
    wire N__5879;
    wire N__5876;
    wire N__5875;
    wire N__5870;
    wire N__5867;
    wire N__5866;
    wire N__5863;
    wire N__5860;
    wire N__5855;
    wire N__5854;
    wire N__5853;
    wire N__5852;
    wire N__5849;
    wire N__5842;
    wire N__5839;
    wire N__5834;
    wire N__5831;
    wire N__5828;
    wire N__5827;
    wire N__5824;
    wire N__5823;
    wire N__5822;
    wire N__5821;
    wire N__5820;
    wire N__5817;
    wire N__5814;
    wire N__5811;
    wire N__5808;
    wire N__5803;
    wire N__5800;
    wire N__5797;
    wire N__5794;
    wire N__5789;
    wire N__5784;
    wire N__5777;
    wire N__5774;
    wire N__5771;
    wire N__5768;
    wire N__5767;
    wire N__5764;
    wire N__5763;
    wire N__5762;
    wire N__5761;
    wire N__5760;
    wire N__5757;
    wire N__5754;
    wire N__5749;
    wire N__5748;
    wire N__5747;
    wire N__5746;
    wire N__5743;
    wire N__5742;
    wire N__5741;
    wire N__5738;
    wire N__5735;
    wire N__5732;
    wire N__5729;
    wire N__5722;
    wire N__5719;
    wire N__5714;
    wire N__5711;
    wire N__5702;
    wire N__5697;
    wire N__5694;
    wire N__5689;
    wire N__5684;
    wire N__5683;
    wire N__5682;
    wire N__5681;
    wire N__5680;
    wire N__5679;
    wire N__5676;
    wire N__5675;
    wire N__5674;
    wire N__5673;
    wire N__5668;
    wire N__5665;
    wire N__5662;
    wire N__5659;
    wire N__5656;
    wire N__5653;
    wire N__5648;
    wire N__5645;
    wire N__5644;
    wire N__5643;
    wire N__5640;
    wire N__5637;
    wire N__5634;
    wire N__5631;
    wire N__5626;
    wire N__5623;
    wire N__5618;
    wire N__5611;
    wire N__5602;
    wire N__5597;
    wire N__5594;
    wire N__5591;
    wire N__5590;
    wire N__5587;
    wire N__5584;
    wire N__5581;
    wire N__5578;
    wire N__5575;
    wire N__5572;
    wire N__5567;
    wire N__5564;
    wire N__5563;
    wire N__5562;
    wire N__5561;
    wire N__5558;
    wire N__5555;
    wire N__5550;
    wire N__5549;
    wire N__5548;
    wire N__5547;
    wire N__5546;
    wire N__5545;
    wire N__5542;
    wire N__5539;
    wire N__5536;
    wire N__5531;
    wire N__5526;
    wire N__5523;
    wire N__5510;
    wire N__5507;
    wire N__5504;
    wire N__5501;
    wire N__5500;
    wire N__5499;
    wire N__5498;
    wire N__5497;
    wire N__5496;
    wire N__5495;
    wire N__5494;
    wire N__5491;
    wire N__5488;
    wire N__5483;
    wire N__5478;
    wire N__5475;
    wire N__5472;
    wire N__5469;
    wire N__5456;
    wire N__5455;
    wire N__5452;
    wire N__5449;
    wire N__5448;
    wire N__5447;
    wire N__5446;
    wire N__5445;
    wire N__5444;
    wire N__5443;
    wire N__5440;
    wire N__5437;
    wire N__5430;
    wire N__5427;
    wire N__5422;
    wire N__5419;
    wire N__5408;
    wire N__5407;
    wire N__5406;
    wire N__5405;
    wire N__5402;
    wire N__5399;
    wire N__5398;
    wire N__5397;
    wire N__5394;
    wire N__5391;
    wire N__5388;
    wire N__5385;
    wire N__5380;
    wire N__5377;
    wire N__5366;
    wire N__5365;
    wire N__5364;
    wire N__5363;
    wire N__5362;
    wire N__5359;
    wire N__5354;
    wire N__5351;
    wire N__5350;
    wire N__5347;
    wire N__5342;
    wire N__5339;
    wire N__5334;
    wire N__5327;
    wire N__5326;
    wire N__5325;
    wire N__5322;
    wire N__5317;
    wire N__5312;
    wire N__5311;
    wire N__5310;
    wire N__5309;
    wire N__5306;
    wire N__5303;
    wire N__5300;
    wire N__5299;
    wire N__5296;
    wire N__5295;
    wire N__5292;
    wire N__5291;
    wire N__5290;
    wire N__5285;
    wire N__5282;
    wire N__5281;
    wire N__5278;
    wire N__5275;
    wire N__5272;
    wire N__5267;
    wire N__5264;
    wire N__5259;
    wire N__5246;
    wire N__5243;
    wire N__5240;
    wire N__5237;
    wire N__5234;
    wire N__5231;
    wire N__5228;
    wire N__5225;
    wire N__5222;
    wire N__5219;
    wire N__5218;
    wire N__5217;
    wire N__5216;
    wire N__5213;
    wire N__5210;
    wire N__5207;
    wire N__5204;
    wire N__5203;
    wire N__5202;
    wire N__5197;
    wire N__5192;
    wire N__5189;
    wire N__5188;
    wire N__5185;
    wire N__5182;
    wire N__5179;
    wire N__5176;
    wire N__5173;
    wire N__5170;
    wire N__5165;
    wire N__5156;
    wire N__5155;
    wire N__5154;
    wire N__5151;
    wire N__5148;
    wire N__5147;
    wire N__5144;
    wire N__5139;
    wire N__5138;
    wire N__5135;
    wire N__5134;
    wire N__5133;
    wire N__5130;
    wire N__5127;
    wire N__5120;
    wire N__5117;
    wire N__5108;
    wire N__5105;
    wire N__5102;
    wire N__5099;
    wire N__5096;
    wire N__5093;
    wire N__5092;
    wire N__5089;
    wire N__5088;
    wire N__5085;
    wire N__5082;
    wire N__5079;
    wire N__5078;
    wire N__5075;
    wire N__5070;
    wire N__5067;
    wire N__5060;
    wire N__5057;
    wire N__5054;
    wire N__5051;
    wire N__5048;
    wire N__5045;
    wire N__5042;
    wire N__5039;
    wire N__5036;
    wire N__5033;
    wire N__5030;
    wire N__5029;
    wire N__5026;
    wire N__5023;
    wire N__5020;
    wire N__5015;
    wire N__5014;
    wire N__5009;
    wire N__5006;
    wire N__5005;
    wire N__5004;
    wire N__5003;
    wire N__5002;
    wire N__4999;
    wire N__4992;
    wire N__4989;
    wire N__4982;
    wire N__4981;
    wire N__4980;
    wire N__4977;
    wire N__4972;
    wire N__4969;
    wire N__4966;
    wire N__4965;
    wire N__4964;
    wire N__4963;
    wire N__4958;
    wire N__4953;
    wire N__4950;
    wire N__4943;
    wire N__4940;
    wire N__4937;
    wire N__4934;
    wire N__4931;
    wire N__4928;
    wire N__4925;
    wire N__4922;
    wire N__4919;
    wire N__4916;
    wire N__4913;
    wire N__4910;
    wire N__4907;
    wire N__4904;
    wire N__4901;
    wire N__4898;
    wire N__4897;
    wire N__4894;
    wire N__4891;
    wire N__4890;
    wire N__4889;
    wire N__4884;
    wire N__4879;
    wire N__4874;
    wire N__4871;
    wire N__4868;
    wire N__4865;
    wire N__4862;
    wire N__4859;
    wire N__4856;
    wire N__4853;
    wire N__4850;
    wire N__4847;
    wire N__4844;
    wire N__4841;
    wire N__4838;
    wire N__4837;
    wire N__4834;
    wire N__4833;
    wire N__4832;
    wire N__4829;
    wire N__4826;
    wire N__4823;
    wire N__4820;
    wire N__4817;
    wire N__4808;
    wire N__4807;
    wire N__4806;
    wire N__4805;
    wire N__4804;
    wire N__4803;
    wire N__4802;
    wire N__4801;
    wire N__4800;
    wire N__4799;
    wire N__4798;
    wire N__4797;
    wire N__4796;
    wire N__4795;
    wire N__4794;
    wire N__4793;
    wire N__4792;
    wire N__4791;
    wire N__4790;
    wire N__4789;
    wire N__4788;
    wire N__4787;
    wire N__4786;
    wire N__4785;
    wire N__4784;
    wire N__4783;
    wire N__4782;
    wire N__4781;
    wire N__4780;
    wire N__4779;
    wire N__4778;
    wire N__4777;
    wire N__4776;
    wire N__4775;
    wire N__4774;
    wire N__4773;
    wire N__4700;
    wire N__4697;
    wire N__4694;
    wire N__4693;
    wire N__4692;
    wire N__4691;
    wire N__4690;
    wire N__4687;
    wire N__4686;
    wire N__4681;
    wire N__4678;
    wire N__4673;
    wire N__4670;
    wire N__4669;
    wire N__4668;
    wire N__4667;
    wire N__4666;
    wire N__4663;
    wire N__4658;
    wire N__4655;
    wire N__4654;
    wire N__4651;
    wire N__4648;
    wire N__4645;
    wire N__4644;
    wire N__4641;
    wire N__4640;
    wire N__4639;
    wire N__4632;
    wire N__4629;
    wire N__4626;
    wire N__4623;
    wire N__4620;
    wire N__4615;
    wire N__4610;
    wire N__4607;
    wire N__4604;
    wire N__4589;
    wire N__4588;
    wire N__4587;
    wire N__4584;
    wire N__4581;
    wire N__4580;
    wire N__4579;
    wire N__4578;
    wire N__4577;
    wire N__4574;
    wire N__4571;
    wire N__4568;
    wire N__4563;
    wire N__4558;
    wire N__4555;
    wire N__4548;
    wire N__4547;
    wire N__4544;
    wire N__4543;
    wire N__4542;
    wire N__4541;
    wire N__4540;
    wire N__4539;
    wire N__4536;
    wire N__4533;
    wire N__4530;
    wire N__4527;
    wire N__4522;
    wire N__4515;
    wire N__4502;
    wire N__4501;
    wire N__4498;
    wire N__4497;
    wire N__4494;
    wire N__4493;
    wire N__4492;
    wire N__4489;
    wire N__4486;
    wire N__4485;
    wire N__4482;
    wire N__4479;
    wire N__4476;
    wire N__4473;
    wire N__4470;
    wire N__4467;
    wire N__4462;
    wire N__4459;
    wire N__4458;
    wire N__4457;
    wire N__4454;
    wire N__4447;
    wire N__4444;
    wire N__4439;
    wire N__4430;
    wire N__4427;
    wire N__4424;
    wire N__4421;
    wire N__4418;
    wire N__4417;
    wire N__4414;
    wire N__4413;
    wire N__4412;
    wire N__4411;
    wire N__4408;
    wire N__4405;
    wire N__4402;
    wire N__4397;
    wire N__4388;
    wire N__4387;
    wire N__4384;
    wire N__4383;
    wire N__4380;
    wire N__4377;
    wire N__4374;
    wire N__4369;
    wire N__4366;
    wire N__4363;
    wire N__4358;
    wire N__4355;
    wire N__4352;
    wire N__4351;
    wire N__4348;
    wire N__4345;
    wire N__4340;
    wire N__4337;
    wire N__4334;
    wire N__4331;
    wire N__4328;
    wire N__4325;
    wire N__4322;
    wire N__4319;
    wire N__4316;
    wire N__4313;
    wire N__4310;
    wire N__4309;
    wire N__4308;
    wire N__4305;
    wire N__4302;
    wire N__4299;
    wire N__4292;
    wire N__4289;
    wire N__4286;
    wire N__4283;
    wire N__4280;
    wire N__4277;
    wire N__4274;
    wire N__4273;
    wire N__4272;
    wire N__4271;
    wire N__4268;
    wire N__4267;
    wire N__4264;
    wire N__4259;
    wire N__4256;
    wire N__4253;
    wire N__4252;
    wire N__4251;
    wire N__4250;
    wire N__4249;
    wire N__4248;
    wire N__4243;
    wire N__4238;
    wire N__4233;
    wire N__4228;
    wire N__4225;
    wire N__4214;
    wire N__4213;
    wire N__4210;
    wire N__4207;
    wire N__4206;
    wire N__4205;
    wire N__4204;
    wire N__4203;
    wire N__4198;
    wire N__4195;
    wire N__4194;
    wire N__4191;
    wire N__4188;
    wire N__4185;
    wire N__4184;
    wire N__4183;
    wire N__4180;
    wire N__4179;
    wire N__4176;
    wire N__4173;
    wire N__4166;
    wire N__4161;
    wire N__4158;
    wire N__4155;
    wire N__4150;
    wire N__4147;
    wire N__4136;
    wire N__4135;
    wire N__4132;
    wire N__4129;
    wire N__4126;
    wire N__4121;
    wire N__4118;
    wire N__4117;
    wire N__4112;
    wire N__4109;
    wire N__4106;
    wire N__4103;
    wire N__4100;
    wire N__4097;
    wire N__4094;
    wire N__4091;
    wire N__4088;
    wire N__4085;
    wire N__4082;
    wire N__4079;
    wire N__4076;
    wire N__4073;
    wire N__4070;
    wire N__4067;
    wire N__4064;
    wire N__4061;
    wire N__4058;
    wire N__4055;
    wire N__4052;
    wire N__4049;
    wire N__4046;
    wire N__4043;
    wire N__4040;
    wire N__4037;
    wire N__4034;
    wire N__4031;
    wire N__4028;
    wire N__4025;
    wire N__4022;
    wire N__4019;
    wire N__4016;
    wire N__4013;
    wire N__4010;
    wire N__4009;
    wire N__4006;
    wire N__4003;
    wire N__4000;
    wire N__3997;
    wire N__3992;
    wire N__3989;
    wire N__3986;
    wire N__3985;
    wire N__3982;
    wire N__3979;
    wire N__3976;
    wire N__3971;
    wire N__3968;
    wire N__3967;
    wire N__3966;
    wire N__3965;
    wire N__3964;
    wire N__3963;
    wire N__3960;
    wire N__3955;
    wire N__3952;
    wire N__3949;
    wire N__3946;
    wire N__3943;
    wire N__3940;
    wire N__3937;
    wire N__3926;
    wire N__3925;
    wire N__3922;
    wire N__3919;
    wire N__3916;
    wire N__3913;
    wire N__3912;
    wire N__3909;
    wire N__3906;
    wire N__3903;
    wire N__3900;
    wire N__3897;
    wire N__3890;
    wire N__3889;
    wire N__3888;
    wire N__3885;
    wire N__3882;
    wire N__3879;
    wire N__3876;
    wire N__3875;
    wire N__3872;
    wire N__3869;
    wire N__3866;
    wire N__3863;
    wire N__3860;
    wire N__3857;
    wire N__3848;
    wire N__3845;
    wire N__3842;
    wire N__3839;
    wire N__3836;
    wire N__3833;
    wire N__3830;
    wire N__3827;
    wire N__3824;
    wire N__3821;
    wire N__3820;
    wire N__3817;
    wire N__3814;
    wire N__3809;
    wire N__3806;
    wire N__3803;
    wire N__3800;
    wire N__3797;
    wire N__3794;
    wire N__3791;
    wire N__3788;
    wire N__3785;
    wire N__3782;
    wire N__3779;
    wire N__3776;
    wire N__3773;
    wire N__3770;
    wire N__3769;
    wire N__3766;
    wire N__3763;
    wire N__3760;
    wire N__3757;
    wire N__3752;
    wire N__3749;
    wire N__3746;
    wire N__3743;
    wire N__3740;
    wire N__3737;
    wire N__3734;
    wire N__3731;
    wire N__3728;
    wire N__3725;
    wire N__3722;
    wire N__3719;
    wire N__3718;
    wire N__3715;
    wire N__3712;
    wire N__3711;
    wire N__3708;
    wire N__3705;
    wire N__3704;
    wire N__3701;
    wire N__3700;
    wire N__3695;
    wire N__3692;
    wire N__3689;
    wire N__3686;
    wire N__3681;
    wire N__3678;
    wire N__3671;
    wire N__3670;
    wire N__3667;
    wire N__3666;
    wire N__3663;
    wire N__3662;
    wire N__3659;
    wire N__3656;
    wire N__3653;
    wire N__3650;
    wire N__3645;
    wire N__3644;
    wire N__3643;
    wire N__3636;
    wire N__3631;
    wire N__3626;
    wire N__3623;
    wire N__3622;
    wire N__3619;
    wire N__3616;
    wire N__3611;
    wire N__3608;
    wire N__3605;
    wire N__3602;
    wire N__3599;
    wire N__3598;
    wire N__3593;
    wire N__3590;
    wire N__3587;
    wire N__3584;
    wire N__3581;
    wire N__3578;
    wire N__3575;
    wire N__3572;
    wire N__3569;
    wire N__3566;
    wire N__3563;
    wire N__3560;
    wire N__3557;
    wire N__3554;
    wire N__3551;
    wire N__3548;
    wire N__3547;
    wire N__3546;
    wire N__3545;
    wire N__3542;
    wire N__3541;
    wire N__3538;
    wire N__3537;
    wire N__3534;
    wire N__3527;
    wire N__3524;
    wire N__3523;
    wire N__3520;
    wire N__3517;
    wire N__3516;
    wire N__3515;
    wire N__3514;
    wire N__3511;
    wire N__3508;
    wire N__3503;
    wire N__3500;
    wire N__3493;
    wire N__3486;
    wire N__3479;
    wire N__3476;
    wire N__3473;
    wire N__3470;
    wire N__3467;
    wire N__3464;
    wire N__3461;
    wire N__3458;
    wire N__3455;
    wire N__3452;
    wire N__3449;
    wire N__3446;
    wire N__3443;
    wire N__3440;
    wire N__3437;
    wire N__3434;
    wire N__3433;
    wire N__3432;
    wire N__3429;
    wire N__3428;
    wire N__3425;
    wire N__3424;
    wire N__3421;
    wire N__3418;
    wire N__3413;
    wire N__3410;
    wire N__3409;
    wire N__3406;
    wire N__3401;
    wire N__3398;
    wire N__3395;
    wire N__3386;
    wire N__3383;
    wire N__3380;
    wire N__3377;
    wire N__3376;
    wire N__3375;
    wire N__3374;
    wire N__3371;
    wire N__3366;
    wire N__3363;
    wire N__3356;
    wire N__3355;
    wire N__3352;
    wire N__3351;
    wire N__3348;
    wire N__3345;
    wire N__3340;
    wire N__3335;
    wire N__3332;
    wire N__3329;
    wire N__3328;
    wire N__3327;
    wire N__3324;
    wire N__3319;
    wire N__3314;
    wire N__3311;
    wire N__3308;
    wire N__3305;
    wire N__3302;
    wire N__3301;
    wire N__3298;
    wire N__3297;
    wire N__3296;
    wire N__3295;
    wire N__3292;
    wire N__3289;
    wire N__3286;
    wire N__3281;
    wire N__3272;
    wire N__3269;
    wire N__3268;
    wire N__3267;
    wire N__3266;
    wire N__3265;
    wire N__3262;
    wire N__3255;
    wire N__3252;
    wire N__3245;
    wire N__3242;
    wire N__3239;
    wire N__3236;
    wire N__3233;
    wire N__3230;
    wire N__3227;
    wire N__3224;
    wire N__3221;
    wire N__3218;
    wire N__3215;
    wire N__3212;
    wire N__3211;
    wire N__3210;
    wire N__3207;
    wire N__3202;
    wire N__3197;
    wire N__3194;
    wire N__3191;
    wire N__3188;
    wire N__3185;
    wire N__3184;
    wire N__3183;
    wire N__3182;
    wire N__3181;
    wire N__3180;
    wire N__3177;
    wire N__3172;
    wire N__3167;
    wire N__3164;
    wire N__3155;
    wire N__3154;
    wire N__3153;
    wire N__3152;
    wire N__3151;
    wire N__3148;
    wire N__3145;
    wire N__3140;
    wire N__3137;
    wire N__3132;
    wire N__3127;
    wire N__3124;
    wire N__3119;
    wire N__3116;
    wire N__3113;
    wire N__3110;
    wire N__3107;
    wire N__3106;
    wire N__3103;
    wire N__3100;
    wire N__3097;
    wire N__3092;
    wire N__3089;
    wire N__3086;
    wire N__3083;
    wire N__3080;
    wire N__3077;
    wire N__3074;
    wire N__3071;
    wire N__3068;
    wire N__3065;
    wire N__3062;
    wire N__3059;
    wire N__3056;
    wire N__3053;
    wire N__3050;
    wire N__3047;
    wire N__3044;
    wire N__3041;
    wire N__3038;
    wire N__3035;
    wire N__3032;
    wire N__3029;
    wire N__3026;
    wire N__3023;
    wire N__3020;
    wire N__3017;
    wire N__3014;
    wire N__3011;
    wire N__3008;
    wire N__3007;
    wire N__3002;
    wire N__2999;
    wire N__2998;
    wire N__2995;
    wire N__2992;
    wire N__2989;
    wire N__2984;
    wire N__2981;
    wire N__2978;
    wire N__2975;
    wire N__2972;
    wire N__2969;
    wire N__2966;
    wire N__2963;
    wire N__2960;
    wire N__2957;
    wire N__2954;
    wire N__2951;
    wire N__2948;
    wire N__2945;
    wire N__2942;
    wire N__2939;
    wire N__2936;
    wire N__2933;
    wire N__2930;
    wire N__2927;
    wire N__2924;
    wire N__2921;
    wire N__2918;
    wire N__2915;
    wire N__2912;
    wire N__2909;
    wire N__2906;
    wire N__2903;
    wire N__2900;
    wire N__2897;
    wire N__2894;
    wire N__2891;
    wire N__2888;
    wire N__2885;
    wire N__2882;
    wire N__2879;
    wire N__2876;
    wire N__2873;
    wire N__2870;
    wire N__2867;
    wire N__2864;
    wire N__2861;
    wire N__2858;
    wire N__2855;
    wire N__2852;
    wire N__2849;
    wire GNDG0;
    wire VCCG0;
    wire \INVseq.counter.T_0_2_rep1C_net ;
    wire clk_c;
    wire buf_clk_1;
    wire \pc.N_21_0_cascade_ ;
    wire seq_D_6_cascade_;
    wire \pc.G_12_i_a3_1 ;
    wire \pc.program_counter_m_3_cascade_ ;
    wire \pc.tbuf.gZ0Z3 ;
    wire \pc.tbuf.g0Z0Z_3_cascade_ ;
    wire bus_3_cascade_;
    wire \INVAR.ff4.qC_net ;
    wire seq_MAR_LD_1_0;
    wire \pc.program_counter_m_3 ;
    wire \seq.DZ0Z_0_cascade_ ;
    wire seq_un1_IR_OE_4_1_cascade_;
    wire \pc.program_counter_RNO_5Z0Z_0 ;
    wire \seq.un17_IR_OE_cascade_ ;
    wire seq_PC_LD_0_0_cascade_;
    wire \seq.D_6_x ;
    wire \INVIR.ff5.q_0_rep1C_net ;
    wire bus_6_cascade_;
    wire N_5_0_cascade_;
    wire \INVIR.ff7.q_ret_1C_net ;
    wire \INVIR.ff5.q_0_nerC_net ;
    wire \INVseq.counter.T_4C_net ;
    wire mem_data_2_7_0__g1;
    wire \pc.program_counter_m_0_2_cascade_ ;
    wire AR_out_2;
    wire \INVAR.ff3.qC_net ;
    wire AR_out_0;
    wire mem_data_2_7_0__N_7_0;
    wire \pc.program_counter_m_0_0 ;
    wire \pc.out_1_2_iv_0_cascade_ ;
    wire \pc.tbuf.g0Z0Z_1_cascade_ ;
    wire bus_0;
    wire mem_data_2_7_0__N_14_0;
    wire \ALU_main.N_48_cascade_ ;
    wire alu_out_m_7_cascade_;
    wire acc_out_m_7_cascade_;
    wire out_c_7;
    wire \INVout_reg.ff8.qC_net ;
    wire \pc.out_1_2_iv_0 ;
    wire \pc.program_counter_RNO_7Z0Z_0_cascade_ ;
    wire \pc.program_counter_RNO_3Z0Z_0 ;
    wire \pc.program_counter_RNO_8Z0Z_0 ;
    wire \INVmar.ff1.q_nerC_net ;
    wire ROM_OE_cascade_;
    wire \pc.program_counter_m_2 ;
    wire \pc.out_1_0_iv_0 ;
    wire \pc.G_10_0_a11_2_1_cascade_ ;
    wire \pc.N_23 ;
    wire \pc.program_counter_RNO_6Z0Z_2_cascade_ ;
    wire \pc.G_10_0_a11_5_2 ;
    wire \seq.S1_1Z0Z_0_cascade_ ;
    wire seq_S1_0_cascade_;
    wire \pc.N_16 ;
    wire bus_6;
    wire ir_out_fast_4;
    wire \seq.counter.T_RNI0T6TZ0Z_4_cascade_ ;
    wire ir_out_7_rep1;
    wire \INVIR.ff7.q_0_fastC_net ;
    wire seq_T_2_rep1;
    wire \seq.D_1_0_x_cascade_ ;
    wire \INVIR.ff6.q_ret_1C_net ;
    wire \seq.B_LD_0_2_tz_cascade_ ;
    wire \seq.counter.T_RNIR83I4_0Z0Z_3 ;
    wire IR_ff6_q_0_fast;
    wire IR_ff7_q_ret_1_fast;
    wire \seq.counter.T_0_fast_RNIP4D21Z0Z_2_cascade_ ;
    wire T_0_fast_RNILB791_2_cascade_;
    wire \pc.G_12_i_0 ;
    wire \seq.counter.T_0_fast_RNIG89VZ0Z_2_cascade_ ;
    wire ir_out_fast_7;
    wire \INVseq.counter.T_0_fast_2C_net ;
    wire \seq.S0_0_i_N_3LZ0Z3 ;
    wire ir_out_i_2_6;
    wire \INVIR.ff7.q_0_nerC_net ;
    wire \seq.counter.T_fast_2 ;
    wire seq_un1_IR_OE_4_1;
    wire g0_0_1_cascade_;
    wire \seq.counter.un7_ACC_LD_0 ;
    wire \seq.un1_ALU_en_0Z0Z_1 ;
    wire \seq.counter.un7_ACC_LD_0_cascade_ ;
    wire IR_OE_2_cascade_;
    wire bus_2;
    wire \seq.g2Z0Z_0 ;
    wire IR_OE_1_cascade_;
    wire \pc.un1_inc_0 ;
    wire \pc.G_12_i_a3_2_3 ;
    wire \pc.G_12_i_a3_2_1 ;
    wire \seq.counter.T8_1_cascade_ ;
    wire \pc.g1_0 ;
    wire \pc.N_188_0 ;
    wire seq_T_0;
    wire \INVseq.counter.T_0C_net ;
    wire N_30;
    wire \pc.G_10_0_1_0_cascade_ ;
    wire \pc.G_10_0_sx ;
    wire \pc.G_10_0_5_1 ;
    wire ALU_main_N_43_0;
    wire \pc.program_counterZ0Z_2 ;
    wire \pc.program_counterZ0Z_0 ;
    wire seq_S0_0_i;
    wire bfn_4_12_0_;
    wire \ALU_main.un1_A_cry_0_c_THRU_CO ;
    wire \ALU_main.un1_A_cry_0 ;
    wire \ALU_main.un1_A_axb_2_l_ofxZ0 ;
    wire un1_A_cry_1_c_RNITKPO2;
    wire \ALU_main.un1_A_cry_1 ;
    wire \ALU_main.un1_A_cry_2 ;
    wire \ALU_main.un1_A_cry_3 ;
    wire \ALU_main.un1_A_cry_4 ;
    wire \ALU_main.un1_A_cry_5 ;
    wire \ALU_main.un1_A_cry_6 ;
    wire bfn_4_13_0_;
    wire \ALU_main.un1_A_cry_6_c_RNIP89EZ0Z2 ;
    wire \ALU_main.un1_A_cry_5_c_RNIDLAPZ0Z2 ;
    wire ALU_main_N_44_0_cascade_;
    wire un1_A_cry_2_c_RNI1TTO2;
    wire \pc.N_10_i ;
    wire \pc.G_10_0_1_1 ;
    wire \pc.G_10_0_1 ;
    wire ALU_main_N_44_1;
    wire \pc.un1_inc_0_0 ;
    wire \pc.out_1_iv_1_1 ;
    wire mem_data_2_7_0__N_16_0;
    wire \pc.g0_rn_1 ;
    wire \pc.g0_sn_cascade_ ;
    wire alu_out_m_0_3;
    wire \pc.program_counterZ0Z_3 ;
    wire seq_un1_AR_OE_0_0;
    wire ir_out_6;
    wire \AR.ff4.AR_out_3 ;
    wire ir_out_3;
    wire \pc.tbuf.g0_0_1_0 ;
    wire AR_out_m_3_cascade_;
    wire \pc.g0_0 ;
    wire ir_out_5;
    wire bus_7;
    wire N_5_0;
    wire N_1_0_cascade_;
    wire seq_un1_HLT_0;
    wire \INVseq.q_ret_1C_net ;
    wire \seq.un1_HLT_1_reti ;
    wire N_2_0;
    wire \seq.un1_HLT_1 ;
    wire \INVseq.q_retC_net ;
    wire bus_1_cascade_;
    wire seq_D_6;
    wire T_0_fast_RNILB791_2;
    wire AR_out_1;
    wire \INVAR.ff2.qC_net ;
    wire \seq.D_3 ;
    wire \seq.counter.ACC_LD_0_0_cascade_ ;
    wire \pc.program_counter_m_0_1 ;
    wire \pc.tbuf.out_1_1_ivZ0Z_0 ;
    wire mem_data_2_7_0__N_11_0_cascade_;
    wire \pc.program_counter_4_rn_2_1 ;
    wire \pc.program_counter_4_sn_1 ;
    wire \pc.g0_1_0_cascade_ ;
    wire \pc.program_counterZ0Z_1 ;
    wire buf_clk_1_g;
    wire seq_T_2;
    wire seq_PC_LD_0_0;
    wire seq_MAR_LD_2;
    wire \seq.gZ0Z2 ;
    wire ALU_main_N_42_0_cascade_;
    wire un1_A_cry_0_c_RNIPCLO2;
    wire ALU_main_N_41_0_cascade_;
    wire un1_A_cry_0_s;
    wire \seq.D_4 ;
    wire \seq.DZ0Z_0 ;
    wire \seq.g2Z0Z_1 ;
    wire \ALU_main.un1_A_axb_0_l_ofxZ0 ;
    wire \ALU_main.un1_A_axb_3_l_ofxZ0 ;
    wire \ALU_main.un1_A_cry_4_c_RNI9D6PZ0Z2 ;
    wire \ALU_main.N_46_cascade_ ;
    wire ir_out_i_2_5;
    wire ir_out_4_rep1;
    wire IR_ff7_q_0_fast;
    wire \seq.counter.TZ0Z_4 ;
    wire ir_out_7;
    wire \seq.g0_i_a3_0Z0Z_2_cascade_ ;
    wire \seq.g0_i_a3Z0Z_2 ;
    wire seq_S0_0_cascade_;
    wire \ALU_main.un1_A_axb_5_l_ofxZ0 ;
    wire \seq.counter.TZ0Z_3 ;
    wire \seq.D_2 ;
    wire \seq.B_LD_0_2_tz ;
    wire \seq.D_1 ;
    wire \ALU_main.un1_A_axb_1_l_ofxZ0 ;
    wire \INVb_reg.ff5.qC_net ;
    wire \ALU_main.un1_A_axb_4_l_ofxZ0 ;
    wire \ALU_main.N_47 ;
    wire acc_out_6;
    wire \ALU_main.un1_A_axb_6_l_ofxZ0 ;
    wire acc_out_7;
    wire acc_out_5;
    wire acc_out_3;
    wire \INVacc.ff7.qC_net ;
    wire \ALU_main.un1_A_cry_3_c_RNI552PZ0Z2 ;
    wire seq_un1_ALU_en_0;
    wire seq_S1_0;
    wire alu_out_m_4_cascade_;
    wire bus_4;
    wire bus_4_cascade_;
    wire ir_out_4;
    wire N_4_0;
    wire b_reg_out_4;
    wire seq_S0_0;
    wire \ALU_main.N_45 ;
    wire bus_5;
    wire \INVIR.ff2.q_nerC_net ;
    wire acc_out_0;
    wire acc_out_1;
    wire acc_out_2;
    wire \INVacc.ff1.qC_net ;
    wire seq_ACC_LD_0_i;
    wire \INVmar.ff4.q_nerC_net ;
    wire \mar.MAR_LD_0_0 ;
    wire b_reg_out_5;
    wire acc_out_m_7;
    wire alu_out_m_7;
    wire b_reg_out_7;
    wire b_reg_out_0;
    wire \INVb_reg.ff6.qC_net ;
    wire \mem.i2_mux_cascade_ ;
    wire \pc.N_7 ;
    wire mem_data_2_7_0__N_29_mux_cascade_;
    wire out_c_6;
    wire \INVout_reg.ff7.qC_net ;
    wire mar_out_2;
    wire mar_out_1;
    wire mar_out_3;
    wire mar_out_0;
    wire mem_data_2_7_0__i2_mux_0;
    wire b_reg_out_1;
    wire acc_out_m_6;
    wire alu_out_m_6;
    wire mem_data_2_7_0__N_29_mux;
    wire b_reg_out_6;
    wire \INVb_reg.ff2.qC_net ;
    wire acc_out_m_5;
    wire alu_out_m_5;
    wire m20;
    wire ROM_OE;
    wire out_c_5;
    wire \INVout_reg.ff6.qC_net ;
    wire out_c_2;
    wire out_c_0;
    wire \INVout_reg.ff3.qC_net ;
    wire \pc.tbuf.g0Z0Z_1 ;
    wire IR_OE_0;
    wire alu_out_m_0_0;
    wire ir_out_0;
    wire \INVIR.ff1.q_nerC_net ;
    wire inc;
    wire alu_out_m_0_2;
    wire ir_out_2;
    wire IR_OE_2;
    wire \pc.tbuf.g0_1_1 ;
    wire b_reg_out_2;
    wire \INVb_reg.ff3.qC_net ;
    wire IR_OE_1;
    wire \pc.g0_1_0 ;
    wire ir_out_1;
    wire alu_out_m_0_1;
    wire out_c_1;
    wire alu_out_m_4;
    wire mem_data_2_7_0__i2_mux_i_m;
    wire acc_out_4;
    wire out_c_4;
    wire \INVout_reg.ff2.qC_net ;
    wire b_reg_out_3;
    wire \INVb_reg.ff4.qC_net ;
    wire seq_B_LD_0_i;
    wire \pc.tbuf.g0_0_0 ;
    wire \pc.tbuf.g0Z0Z_3 ;
    wire \pc.tbuf.gZ0Z2 ;
    wire alu_out_m_1_3;
    wire out_c_3;
    wire _gnd_net_;
    wire \INVout_reg.ff4.qC_net ;
    wire OUT_LD;
    wire clr_c_g;

    PRE_IO_GBUF clr_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__9027),
            .GLOBALBUFFEROUTPUT(clr_c_g));
    IO_PAD clr_ibuf_gb_io_iopad (
            .OE(N__9029),
            .DIN(N__9028),
            .DOUT(N__9027),
            .PACKAGEPIN(clr));
    defparam clr_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam clr_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO clr_ibuf_gb_io_preio (
            .PADOEN(N__9029),
            .PADOUT(N__9028),
            .PADIN(N__9027),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD out_obuf_7_iopad (
            .OE(N__9018),
            .DIN(N__9017),
            .DOUT(N__9016),
            .PACKAGEPIN(out[7]));
    defparam out_obuf_7_preio.NEG_TRIGGER=1'b0;
    defparam out_obuf_7_preio.PIN_TYPE=6'b011001;
    PRE_IO out_obuf_7_preio (
            .PADOEN(N__9018),
            .PADOUT(N__9017),
            .PADIN(N__9016),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3047),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam out_obuf_4_iopad.PULLUP=1'b0;
    defparam out_obuf_4_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD out_obuf_4_iopad (
            .OE(N__9009),
            .DIN(N__9008),
            .DOUT(N__9007),
            .PACKAGEPIN(out[4]));
    defparam out_obuf_4_preio.NEG_TRIGGER=1'b0;
    defparam out_obuf_4_preio.PIN_TYPE=6'b011001;
    PRE_IO out_obuf_4_preio (
            .PADOEN(N__9009),
            .PADOUT(N__9008),
            .PADIN(N__9007),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7844),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam out_obuf_3_iopad.PULLUP=1'b0;
    defparam out_obuf_3_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD out_obuf_3_iopad (
            .OE(N__9000),
            .DIN(N__8999),
            .DOUT(N__8998),
            .PACKAGEPIN(out[3]));
    defparam out_obuf_3_preio.NEG_TRIGGER=1'b0;
    defparam out_obuf_3_preio.PIN_TYPE=6'b011001;
    PRE_IO out_obuf_3_preio (
            .PADOEN(N__9000),
            .PADOUT(N__8999),
            .PADIN(N__8998),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7493),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD out_obuf_6_iopad (
            .OE(N__8991),
            .DIN(N__8990),
            .DOUT(N__8989),
            .PACKAGEPIN(out[6]));
    defparam out_obuf_6_preio.NEG_TRIGGER=1'b0;
    defparam out_obuf_6_preio.PIN_TYPE=6'b011001;
    PRE_IO out_obuf_6_preio (
            .PADOEN(N__8991),
            .PADOUT(N__8990),
            .PADIN(N__8989),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__7205),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD out_obuf_5_iopad (
            .OE(N__8982),
            .DIN(N__8981),
            .DOUT(N__8980),
            .PACKAGEPIN(out[5]));
    defparam out_obuf_5_preio.NEG_TRIGGER=1'b0;
    defparam out_obuf_5_preio.PIN_TYPE=6'b011001;
    PRE_IO out_obuf_5_preio (
            .PADOEN(N__8982),
            .PADOUT(N__8981),
            .PADIN(N__8980),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6422),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam out_obuf_0_iopad.PULLUP=1'b0;
    defparam out_obuf_0_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD out_obuf_0_iopad (
            .OE(N__8973),
            .DIN(N__8972),
            .DOUT(N__8971),
            .PACKAGEPIN(out[0]));
    defparam out_obuf_0_preio.NEG_TRIGGER=1'b0;
    defparam out_obuf_0_preio.PIN_TYPE=6'b011001;
    PRE_IO out_obuf_0_preio (
            .PADOEN(N__8973),
            .PADOUT(N__8972),
            .PADIN(N__8971),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6398),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam clk_ibuf_iopad.PULLUP=1'b0;
    defparam clk_ibuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD clk_ibuf_iopad (
            .OE(N__8964),
            .DIN(N__8963),
            .DOUT(N__8962),
            .PACKAGEPIN(clk));
    defparam clk_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam clk_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO clk_ibuf_preio (
            .PADOEN(N__8964),
            .PADOUT(N__8963),
            .PADIN(N__8962),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(clk_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam out_obuf_2_iopad.PULLUP=1'b0;
    defparam out_obuf_2_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD out_obuf_2_iopad (
            .OE(N__8955),
            .DIN(N__8954),
            .DOUT(N__8953),
            .PACKAGEPIN(out[2]));
    defparam out_obuf_2_preio.NEG_TRIGGER=1'b0;
    defparam out_obuf_2_preio.PIN_TYPE=6'b011001;
    PRE_IO out_obuf_2_preio (
            .PADOEN(N__8955),
            .PADOUT(N__8954),
            .PADIN(N__8953),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6407),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam out_obuf_1_iopad.PULLUP=1'b0;
    defparam out_obuf_1_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD out_obuf_1_iopad (
            .OE(N__8946),
            .DIN(N__8945),
            .DOUT(N__8944),
            .PACKAGEPIN(out[1]));
    defparam out_obuf_1_preio.NEG_TRIGGER=1'b0;
    defparam out_obuf_1_preio.PIN_TYPE=6'b011001;
    PRE_IO out_obuf_1_preio (
            .PADOEN(N__8946),
            .PADOUT(N__8945),
            .PADIN(N__8944),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8012),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2290 (
            .O(N__8927),
            .I(N__8923));
    InMux I__2289 (
            .O(N__8926),
            .I(N__8920));
    LocalMux I__2288 (
            .O(N__8923),
            .I(N__8916));
    LocalMux I__2287 (
            .O(N__8920),
            .I(N__8913));
    InMux I__2286 (
            .O(N__8919),
            .I(N__8910));
    Span4Mux_v I__2285 (
            .O(N__8916),
            .I(N__8901));
    Span4Mux_h I__2284 (
            .O(N__8913),
            .I(N__8901));
    LocalMux I__2283 (
            .O(N__8910),
            .I(N__8901));
    InMux I__2282 (
            .O(N__8909),
            .I(N__8898));
    InMux I__2281 (
            .O(N__8908),
            .I(N__8895));
    Span4Mux_h I__2280 (
            .O(N__8901),
            .I(N__8892));
    LocalMux I__2279 (
            .O(N__8898),
            .I(N__8889));
    LocalMux I__2278 (
            .O(N__8895),
            .I(N__8886));
    Odrv4 I__2277 (
            .O(N__8892),
            .I(\pc.tbuf.g0Z0Z_1 ));
    Odrv12 I__2276 (
            .O(N__8889),
            .I(\pc.tbuf.g0Z0Z_1 ));
    Odrv4 I__2275 (
            .O(N__8886),
            .I(\pc.tbuf.g0Z0Z_1 ));
    CascadeMux I__2274 (
            .O(N__8879),
            .I(N__8874));
    CascadeMux I__2273 (
            .O(N__8878),
            .I(N__8870));
    InMux I__2272 (
            .O(N__8877),
            .I(N__8867));
    InMux I__2271 (
            .O(N__8874),
            .I(N__8864));
    InMux I__2270 (
            .O(N__8873),
            .I(N__8861));
    InMux I__2269 (
            .O(N__8870),
            .I(N__8857));
    LocalMux I__2268 (
            .O(N__8867),
            .I(N__8854));
    LocalMux I__2267 (
            .O(N__8864),
            .I(N__8849));
    LocalMux I__2266 (
            .O(N__8861),
            .I(N__8849));
    CascadeMux I__2265 (
            .O(N__8860),
            .I(N__8845));
    LocalMux I__2264 (
            .O(N__8857),
            .I(N__8842));
    Span4Mux_v I__2263 (
            .O(N__8854),
            .I(N__8839));
    Span4Mux_v I__2262 (
            .O(N__8849),
            .I(N__8836));
    InMux I__2261 (
            .O(N__8848),
            .I(N__8833));
    InMux I__2260 (
            .O(N__8845),
            .I(N__8830));
    Span4Mux_s2_h I__2259 (
            .O(N__8842),
            .I(N__8825));
    Span4Mux_s2_h I__2258 (
            .O(N__8839),
            .I(N__8825));
    Odrv4 I__2257 (
            .O(N__8836),
            .I(IR_OE_0));
    LocalMux I__2256 (
            .O(N__8833),
            .I(IR_OE_0));
    LocalMux I__2255 (
            .O(N__8830),
            .I(IR_OE_0));
    Odrv4 I__2254 (
            .O(N__8825),
            .I(IR_OE_0));
    InMux I__2253 (
            .O(N__8816),
            .I(N__8811));
    InMux I__2252 (
            .O(N__8815),
            .I(N__8808));
    InMux I__2251 (
            .O(N__8814),
            .I(N__8804));
    LocalMux I__2250 (
            .O(N__8811),
            .I(N__8799));
    LocalMux I__2249 (
            .O(N__8808),
            .I(N__8799));
    InMux I__2248 (
            .O(N__8807),
            .I(N__8796));
    LocalMux I__2247 (
            .O(N__8804),
            .I(N__8791));
    Span4Mux_v I__2246 (
            .O(N__8799),
            .I(N__8788));
    LocalMux I__2245 (
            .O(N__8796),
            .I(N__8785));
    InMux I__2244 (
            .O(N__8795),
            .I(N__8782));
    InMux I__2243 (
            .O(N__8794),
            .I(N__8779));
    Span4Mux_h I__2242 (
            .O(N__8791),
            .I(N__8776));
    Odrv4 I__2241 (
            .O(N__8788),
            .I(alu_out_m_0_0));
    Odrv4 I__2240 (
            .O(N__8785),
            .I(alu_out_m_0_0));
    LocalMux I__2239 (
            .O(N__8782),
            .I(alu_out_m_0_0));
    LocalMux I__2238 (
            .O(N__8779),
            .I(alu_out_m_0_0));
    Odrv4 I__2237 (
            .O(N__8776),
            .I(alu_out_m_0_0));
    CascadeMux I__2236 (
            .O(N__8765),
            .I(N__8760));
    InMux I__2235 (
            .O(N__8764),
            .I(N__8757));
    InMux I__2234 (
            .O(N__8763),
            .I(N__8752));
    InMux I__2233 (
            .O(N__8760),
            .I(N__8749));
    LocalMux I__2232 (
            .O(N__8757),
            .I(N__8745));
    InMux I__2231 (
            .O(N__8756),
            .I(N__8742));
    CascadeMux I__2230 (
            .O(N__8755),
            .I(N__8739));
    LocalMux I__2229 (
            .O(N__8752),
            .I(N__8736));
    LocalMux I__2228 (
            .O(N__8749),
            .I(N__8733));
    CascadeMux I__2227 (
            .O(N__8748),
            .I(N__8728));
    Span4Mux_v I__2226 (
            .O(N__8745),
            .I(N__8723));
    LocalMux I__2225 (
            .O(N__8742),
            .I(N__8723));
    InMux I__2224 (
            .O(N__8739),
            .I(N__8720));
    Span4Mux_v I__2223 (
            .O(N__8736),
            .I(N__8715));
    Span4Mux_s2_h I__2222 (
            .O(N__8733),
            .I(N__8715));
    InMux I__2221 (
            .O(N__8732),
            .I(N__8712));
    InMux I__2220 (
            .O(N__8731),
            .I(N__8709));
    InMux I__2219 (
            .O(N__8728),
            .I(N__8706));
    Span4Mux_h I__2218 (
            .O(N__8723),
            .I(N__8703));
    LocalMux I__2217 (
            .O(N__8720),
            .I(N__8698));
    Span4Mux_h I__2216 (
            .O(N__8715),
            .I(N__8698));
    LocalMux I__2215 (
            .O(N__8712),
            .I(ir_out_0));
    LocalMux I__2214 (
            .O(N__8709),
            .I(ir_out_0));
    LocalMux I__2213 (
            .O(N__8706),
            .I(ir_out_0));
    Odrv4 I__2212 (
            .O(N__8703),
            .I(ir_out_0));
    Odrv4 I__2211 (
            .O(N__8698),
            .I(ir_out_0));
    CEMux I__2210 (
            .O(N__8687),
            .I(N__8680));
    CascadeMux I__2209 (
            .O(N__8686),
            .I(N__8669));
    CascadeMux I__2208 (
            .O(N__8685),
            .I(N__8656));
    CascadeMux I__2207 (
            .O(N__8684),
            .I(N__8651));
    CEMux I__2206 (
            .O(N__8683),
            .I(N__8648));
    LocalMux I__2205 (
            .O(N__8680),
            .I(N__8645));
    CEMux I__2204 (
            .O(N__8679),
            .I(N__8642));
    CEMux I__2203 (
            .O(N__8678),
            .I(N__8639));
    InMux I__2202 (
            .O(N__8677),
            .I(N__8636));
    InMux I__2201 (
            .O(N__8676),
            .I(N__8633));
    InMux I__2200 (
            .O(N__8675),
            .I(N__8630));
    InMux I__2199 (
            .O(N__8674),
            .I(N__8625));
    InMux I__2198 (
            .O(N__8673),
            .I(N__8625));
    InMux I__2197 (
            .O(N__8672),
            .I(N__8622));
    InMux I__2196 (
            .O(N__8669),
            .I(N__8614));
    InMux I__2195 (
            .O(N__8668),
            .I(N__8614));
    InMux I__2194 (
            .O(N__8667),
            .I(N__8614));
    InMux I__2193 (
            .O(N__8666),
            .I(N__8609));
    InMux I__2192 (
            .O(N__8665),
            .I(N__8609));
    InMux I__2191 (
            .O(N__8664),
            .I(N__8604));
    InMux I__2190 (
            .O(N__8663),
            .I(N__8604));
    InMux I__2189 (
            .O(N__8662),
            .I(N__8601));
    InMux I__2188 (
            .O(N__8661),
            .I(N__8596));
    InMux I__2187 (
            .O(N__8660),
            .I(N__8596));
    InMux I__2186 (
            .O(N__8659),
            .I(N__8587));
    InMux I__2185 (
            .O(N__8656),
            .I(N__8587));
    InMux I__2184 (
            .O(N__8655),
            .I(N__8587));
    InMux I__2183 (
            .O(N__8654),
            .I(N__8587));
    InMux I__2182 (
            .O(N__8651),
            .I(N__8584));
    LocalMux I__2181 (
            .O(N__8648),
            .I(N__8579));
    Sp12to4 I__2180 (
            .O(N__8645),
            .I(N__8579));
    LocalMux I__2179 (
            .O(N__8642),
            .I(N__8576));
    LocalMux I__2178 (
            .O(N__8639),
            .I(N__8573));
    LocalMux I__2177 (
            .O(N__8636),
            .I(N__8568));
    LocalMux I__2176 (
            .O(N__8633),
            .I(N__8568));
    LocalMux I__2175 (
            .O(N__8630),
            .I(N__8563));
    LocalMux I__2174 (
            .O(N__8625),
            .I(N__8563));
    LocalMux I__2173 (
            .O(N__8622),
            .I(N__8560));
    InMux I__2172 (
            .O(N__8621),
            .I(N__8557));
    LocalMux I__2171 (
            .O(N__8614),
            .I(N__8554));
    LocalMux I__2170 (
            .O(N__8609),
            .I(N__8545));
    LocalMux I__2169 (
            .O(N__8604),
            .I(N__8534));
    LocalMux I__2168 (
            .O(N__8601),
            .I(N__8534));
    LocalMux I__2167 (
            .O(N__8596),
            .I(N__8534));
    LocalMux I__2166 (
            .O(N__8587),
            .I(N__8534));
    LocalMux I__2165 (
            .O(N__8584),
            .I(N__8534));
    Span12Mux_s3_h I__2164 (
            .O(N__8579),
            .I(N__8531));
    Span4Mux_h I__2163 (
            .O(N__8576),
            .I(N__8528));
    Span4Mux_h I__2162 (
            .O(N__8573),
            .I(N__8523));
    Span4Mux_s3_v I__2161 (
            .O(N__8568),
            .I(N__8523));
    Span4Mux_s3_v I__2160 (
            .O(N__8563),
            .I(N__8514));
    Span4Mux_s3_h I__2159 (
            .O(N__8560),
            .I(N__8514));
    LocalMux I__2158 (
            .O(N__8557),
            .I(N__8514));
    Span4Mux_s3_h I__2157 (
            .O(N__8554),
            .I(N__8514));
    InMux I__2156 (
            .O(N__8553),
            .I(N__8509));
    InMux I__2155 (
            .O(N__8552),
            .I(N__8509));
    InMux I__2154 (
            .O(N__8551),
            .I(N__8500));
    InMux I__2153 (
            .O(N__8550),
            .I(N__8500));
    InMux I__2152 (
            .O(N__8549),
            .I(N__8500));
    InMux I__2151 (
            .O(N__8548),
            .I(N__8500));
    Span4Mux_v I__2150 (
            .O(N__8545),
            .I(N__8495));
    Span4Mux_v I__2149 (
            .O(N__8534),
            .I(N__8495));
    Odrv12 I__2148 (
            .O(N__8531),
            .I(inc));
    Odrv4 I__2147 (
            .O(N__8528),
            .I(inc));
    Odrv4 I__2146 (
            .O(N__8523),
            .I(inc));
    Odrv4 I__2145 (
            .O(N__8514),
            .I(inc));
    LocalMux I__2144 (
            .O(N__8509),
            .I(inc));
    LocalMux I__2143 (
            .O(N__8500),
            .I(inc));
    Odrv4 I__2142 (
            .O(N__8495),
            .I(inc));
    InMux I__2141 (
            .O(N__8480),
            .I(N__8475));
    InMux I__2140 (
            .O(N__8479),
            .I(N__8472));
    InMux I__2139 (
            .O(N__8478),
            .I(N__8469));
    LocalMux I__2138 (
            .O(N__8475),
            .I(N__8461));
    LocalMux I__2137 (
            .O(N__8472),
            .I(N__8461));
    LocalMux I__2136 (
            .O(N__8469),
            .I(N__8461));
    InMux I__2135 (
            .O(N__8468),
            .I(N__8458));
    Span4Mux_v I__2134 (
            .O(N__8461),
            .I(N__8452));
    LocalMux I__2133 (
            .O(N__8458),
            .I(N__8452));
    InMux I__2132 (
            .O(N__8457),
            .I(N__8449));
    Span4Mux_h I__2131 (
            .O(N__8452),
            .I(N__8443));
    LocalMux I__2130 (
            .O(N__8449),
            .I(N__8443));
    InMux I__2129 (
            .O(N__8448),
            .I(N__8440));
    Odrv4 I__2128 (
            .O(N__8443),
            .I(alu_out_m_0_2));
    LocalMux I__2127 (
            .O(N__8440),
            .I(alu_out_m_0_2));
    InMux I__2126 (
            .O(N__8435),
            .I(N__8431));
    CascadeMux I__2125 (
            .O(N__8434),
            .I(N__8428));
    LocalMux I__2124 (
            .O(N__8431),
            .I(N__8422));
    InMux I__2123 (
            .O(N__8428),
            .I(N__8419));
    InMux I__2122 (
            .O(N__8427),
            .I(N__8416));
    InMux I__2121 (
            .O(N__8426),
            .I(N__8413));
    InMux I__2120 (
            .O(N__8425),
            .I(N__8408));
    Span4Mux_v I__2119 (
            .O(N__8422),
            .I(N__8403));
    LocalMux I__2118 (
            .O(N__8419),
            .I(N__8403));
    LocalMux I__2117 (
            .O(N__8416),
            .I(N__8400));
    LocalMux I__2116 (
            .O(N__8413),
            .I(N__8397));
    InMux I__2115 (
            .O(N__8412),
            .I(N__8394));
    InMux I__2114 (
            .O(N__8411),
            .I(N__8391));
    LocalMux I__2113 (
            .O(N__8408),
            .I(N__8386));
    Span4Mux_v I__2112 (
            .O(N__8403),
            .I(N__8386));
    Odrv4 I__2111 (
            .O(N__8400),
            .I(ir_out_2));
    Odrv12 I__2110 (
            .O(N__8397),
            .I(ir_out_2));
    LocalMux I__2109 (
            .O(N__8394),
            .I(ir_out_2));
    LocalMux I__2108 (
            .O(N__8391),
            .I(ir_out_2));
    Odrv4 I__2107 (
            .O(N__8386),
            .I(ir_out_2));
    CascadeMux I__2106 (
            .O(N__8375),
            .I(N__8370));
    CascadeMux I__2105 (
            .O(N__8374),
            .I(N__8365));
    CascadeMux I__2104 (
            .O(N__8373),
            .I(N__8362));
    InMux I__2103 (
            .O(N__8370),
            .I(N__8359));
    CascadeMux I__2102 (
            .O(N__8369),
            .I(N__8356));
    CascadeMux I__2101 (
            .O(N__8368),
            .I(N__8353));
    InMux I__2100 (
            .O(N__8365),
            .I(N__8350));
    InMux I__2099 (
            .O(N__8362),
            .I(N__8347));
    LocalMux I__2098 (
            .O(N__8359),
            .I(N__8344));
    InMux I__2097 (
            .O(N__8356),
            .I(N__8341));
    InMux I__2096 (
            .O(N__8353),
            .I(N__8338));
    LocalMux I__2095 (
            .O(N__8350),
            .I(N__8335));
    LocalMux I__2094 (
            .O(N__8347),
            .I(N__8332));
    Span4Mux_v I__2093 (
            .O(N__8344),
            .I(N__8325));
    LocalMux I__2092 (
            .O(N__8341),
            .I(N__8325));
    LocalMux I__2091 (
            .O(N__8338),
            .I(N__8325));
    Span4Mux_v I__2090 (
            .O(N__8335),
            .I(N__8322));
    Span4Mux_h I__2089 (
            .O(N__8332),
            .I(N__8319));
    Span4Mux_h I__2088 (
            .O(N__8325),
            .I(N__8316));
    Odrv4 I__2087 (
            .O(N__8322),
            .I(IR_OE_2));
    Odrv4 I__2086 (
            .O(N__8319),
            .I(IR_OE_2));
    Odrv4 I__2085 (
            .O(N__8316),
            .I(IR_OE_2));
    InMux I__2084 (
            .O(N__8309),
            .I(N__8303));
    InMux I__2083 (
            .O(N__8308),
            .I(N__8300));
    InMux I__2082 (
            .O(N__8307),
            .I(N__8297));
    InMux I__2081 (
            .O(N__8306),
            .I(N__8294));
    LocalMux I__2080 (
            .O(N__8303),
            .I(N__8290));
    LocalMux I__2079 (
            .O(N__8300),
            .I(N__8283));
    LocalMux I__2078 (
            .O(N__8297),
            .I(N__8283));
    LocalMux I__2077 (
            .O(N__8294),
            .I(N__8283));
    InMux I__2076 (
            .O(N__8293),
            .I(N__8280));
    Span4Mux_h I__2075 (
            .O(N__8290),
            .I(N__8272));
    Span4Mux_v I__2074 (
            .O(N__8283),
            .I(N__8272));
    LocalMux I__2073 (
            .O(N__8280),
            .I(N__8272));
    InMux I__2072 (
            .O(N__8279),
            .I(N__8269));
    Span4Mux_h I__2071 (
            .O(N__8272),
            .I(N__8266));
    LocalMux I__2070 (
            .O(N__8269),
            .I(N__8263));
    Odrv4 I__2069 (
            .O(N__8266),
            .I(\pc.tbuf.g0_1_1 ));
    Odrv4 I__2068 (
            .O(N__8263),
            .I(\pc.tbuf.g0_1_1 ));
    CascadeMux I__2067 (
            .O(N__8258),
            .I(N__8254));
    InMux I__2066 (
            .O(N__8257),
            .I(N__8246));
    InMux I__2065 (
            .O(N__8254),
            .I(N__8246));
    InMux I__2064 (
            .O(N__8253),
            .I(N__8246));
    LocalMux I__2063 (
            .O(N__8246),
            .I(N__8243));
    Span4Mux_h I__2062 (
            .O(N__8243),
            .I(N__8240));
    Odrv4 I__2061 (
            .O(N__8240),
            .I(b_reg_out_2));
    InMux I__2060 (
            .O(N__8237),
            .I(N__8233));
    InMux I__2059 (
            .O(N__8236),
            .I(N__8230));
    LocalMux I__2058 (
            .O(N__8233),
            .I(N__8223));
    LocalMux I__2057 (
            .O(N__8230),
            .I(N__8223));
    InMux I__2056 (
            .O(N__8229),
            .I(N__8220));
    InMux I__2055 (
            .O(N__8228),
            .I(N__8217));
    Span4Mux_v I__2054 (
            .O(N__8223),
            .I(N__8212));
    LocalMux I__2053 (
            .O(N__8220),
            .I(N__8212));
    LocalMux I__2052 (
            .O(N__8217),
            .I(N__8207));
    Sp12to4 I__2051 (
            .O(N__8212),
            .I(N__8204));
    InMux I__2050 (
            .O(N__8211),
            .I(N__8201));
    InMux I__2049 (
            .O(N__8210),
            .I(N__8198));
    Span12Mux_s7_v I__2048 (
            .O(N__8207),
            .I(N__8193));
    Span12Mux_s8_v I__2047 (
            .O(N__8204),
            .I(N__8193));
    LocalMux I__2046 (
            .O(N__8201),
            .I(N__8188));
    LocalMux I__2045 (
            .O(N__8198),
            .I(N__8188));
    Odrv12 I__2044 (
            .O(N__8193),
            .I(IR_OE_1));
    Odrv4 I__2043 (
            .O(N__8188),
            .I(IR_OE_1));
    InMux I__2042 (
            .O(N__8183),
            .I(N__8179));
    InMux I__2041 (
            .O(N__8182),
            .I(N__8176));
    LocalMux I__2040 (
            .O(N__8179),
            .I(N__8173));
    LocalMux I__2039 (
            .O(N__8176),
            .I(N__8170));
    Span4Mux_v I__2038 (
            .O(N__8173),
            .I(N__8161));
    Span4Mux_h I__2037 (
            .O(N__8170),
            .I(N__8161));
    InMux I__2036 (
            .O(N__8169),
            .I(N__8158));
    InMux I__2035 (
            .O(N__8168),
            .I(N__8155));
    InMux I__2034 (
            .O(N__8167),
            .I(N__8152));
    InMux I__2033 (
            .O(N__8166),
            .I(N__8149));
    Odrv4 I__2032 (
            .O(N__8161),
            .I(\pc.g0_1_0 ));
    LocalMux I__2031 (
            .O(N__8158),
            .I(\pc.g0_1_0 ));
    LocalMux I__2030 (
            .O(N__8155),
            .I(\pc.g0_1_0 ));
    LocalMux I__2029 (
            .O(N__8152),
            .I(\pc.g0_1_0 ));
    LocalMux I__2028 (
            .O(N__8149),
            .I(\pc.g0_1_0 ));
    CascadeMux I__2027 (
            .O(N__8138),
            .I(N__8134));
    CascadeMux I__2026 (
            .O(N__8137),
            .I(N__8131));
    InMux I__2025 (
            .O(N__8134),
            .I(N__8126));
    InMux I__2024 (
            .O(N__8131),
            .I(N__8123));
    CascadeMux I__2023 (
            .O(N__8130),
            .I(N__8118));
    CascadeMux I__2022 (
            .O(N__8129),
            .I(N__8115));
    LocalMux I__2021 (
            .O(N__8126),
            .I(N__8109));
    LocalMux I__2020 (
            .O(N__8123),
            .I(N__8109));
    CascadeMux I__2019 (
            .O(N__8122),
            .I(N__8106));
    CascadeMux I__2018 (
            .O(N__8121),
            .I(N__8103));
    InMux I__2017 (
            .O(N__8118),
            .I(N__8100));
    InMux I__2016 (
            .O(N__8115),
            .I(N__8097));
    InMux I__2015 (
            .O(N__8114),
            .I(N__8094));
    Span4Mux_v I__2014 (
            .O(N__8109),
            .I(N__8091));
    InMux I__2013 (
            .O(N__8106),
            .I(N__8088));
    InMux I__2012 (
            .O(N__8103),
            .I(N__8085));
    LocalMux I__2011 (
            .O(N__8100),
            .I(N__8080));
    LocalMux I__2010 (
            .O(N__8097),
            .I(N__8080));
    LocalMux I__2009 (
            .O(N__8094),
            .I(N__8077));
    Odrv4 I__2008 (
            .O(N__8091),
            .I(ir_out_1));
    LocalMux I__2007 (
            .O(N__8088),
            .I(ir_out_1));
    LocalMux I__2006 (
            .O(N__8085),
            .I(ir_out_1));
    Odrv4 I__2005 (
            .O(N__8080),
            .I(ir_out_1));
    Odrv12 I__2004 (
            .O(N__8077),
            .I(ir_out_1));
    InMux I__2003 (
            .O(N__8066),
            .I(N__8061));
    InMux I__2002 (
            .O(N__8065),
            .I(N__8057));
    InMux I__2001 (
            .O(N__8064),
            .I(N__8054));
    LocalMux I__2000 (
            .O(N__8061),
            .I(N__8049));
    InMux I__1999 (
            .O(N__8060),
            .I(N__8046));
    LocalMux I__1998 (
            .O(N__8057),
            .I(N__8042));
    LocalMux I__1997 (
            .O(N__8054),
            .I(N__8039));
    InMux I__1996 (
            .O(N__8053),
            .I(N__8036));
    InMux I__1995 (
            .O(N__8052),
            .I(N__8033));
    Span4Mux_h I__1994 (
            .O(N__8049),
            .I(N__8028));
    LocalMux I__1993 (
            .O(N__8046),
            .I(N__8028));
    InMux I__1992 (
            .O(N__8045),
            .I(N__8025));
    Odrv4 I__1991 (
            .O(N__8042),
            .I(alu_out_m_0_1));
    Odrv4 I__1990 (
            .O(N__8039),
            .I(alu_out_m_0_1));
    LocalMux I__1989 (
            .O(N__8036),
            .I(alu_out_m_0_1));
    LocalMux I__1988 (
            .O(N__8033),
            .I(alu_out_m_0_1));
    Odrv4 I__1987 (
            .O(N__8028),
            .I(alu_out_m_0_1));
    LocalMux I__1986 (
            .O(N__8025),
            .I(alu_out_m_0_1));
    IoInMux I__1985 (
            .O(N__8012),
            .I(N__8009));
    LocalMux I__1984 (
            .O(N__8009),
            .I(N__8006));
    Odrv12 I__1983 (
            .O(N__8006),
            .I(out_c_1));
    InMux I__1982 (
            .O(N__8003),
            .I(N__7999));
    InMux I__1981 (
            .O(N__8002),
            .I(N__7996));
    LocalMux I__1980 (
            .O(N__7999),
            .I(N__7991));
    LocalMux I__1979 (
            .O(N__7996),
            .I(N__7988));
    InMux I__1978 (
            .O(N__7995),
            .I(N__7985));
    InMux I__1977 (
            .O(N__7994),
            .I(N__7982));
    Span4Mux_v I__1976 (
            .O(N__7991),
            .I(N__7977));
    Span4Mux_h I__1975 (
            .O(N__7988),
            .I(N__7977));
    LocalMux I__1974 (
            .O(N__7985),
            .I(N__7974));
    LocalMux I__1973 (
            .O(N__7982),
            .I(N__7971));
    Odrv4 I__1972 (
            .O(N__7977),
            .I(alu_out_m_4));
    Odrv12 I__1971 (
            .O(N__7974),
            .I(alu_out_m_4));
    Odrv4 I__1970 (
            .O(N__7971),
            .I(alu_out_m_4));
    InMux I__1969 (
            .O(N__7964),
            .I(N__7961));
    LocalMux I__1968 (
            .O(N__7961),
            .I(N__7956));
    InMux I__1967 (
            .O(N__7960),
            .I(N__7953));
    InMux I__1966 (
            .O(N__7959),
            .I(N__7948));
    Span12Mux_s3_v I__1965 (
            .O(N__7956),
            .I(N__7945));
    LocalMux I__1964 (
            .O(N__7953),
            .I(N__7942));
    InMux I__1963 (
            .O(N__7952),
            .I(N__7939));
    InMux I__1962 (
            .O(N__7951),
            .I(N__7936));
    LocalMux I__1961 (
            .O(N__7948),
            .I(N__7933));
    Odrv12 I__1960 (
            .O(N__7945),
            .I(mem_data_2_7_0__i2_mux_i_m));
    Odrv4 I__1959 (
            .O(N__7942),
            .I(mem_data_2_7_0__i2_mux_i_m));
    LocalMux I__1958 (
            .O(N__7939),
            .I(mem_data_2_7_0__i2_mux_i_m));
    LocalMux I__1957 (
            .O(N__7936),
            .I(mem_data_2_7_0__i2_mux_i_m));
    Odrv4 I__1956 (
            .O(N__7933),
            .I(mem_data_2_7_0__i2_mux_i_m));
    CascadeMux I__1955 (
            .O(N__7922),
            .I(N__7919));
    InMux I__1954 (
            .O(N__7919),
            .I(N__7916));
    LocalMux I__1953 (
            .O(N__7916),
            .I(N__7911));
    CascadeMux I__1952 (
            .O(N__7915),
            .I(N__7905));
    CascadeMux I__1951 (
            .O(N__7914),
            .I(N__7900));
    Span4Mux_s2_v I__1950 (
            .O(N__7911),
            .I(N__7897));
    InMux I__1949 (
            .O(N__7910),
            .I(N__7892));
    InMux I__1948 (
            .O(N__7909),
            .I(N__7892));
    CascadeMux I__1947 (
            .O(N__7908),
            .I(N__7889));
    InMux I__1946 (
            .O(N__7905),
            .I(N__7886));
    CascadeMux I__1945 (
            .O(N__7904),
            .I(N__7883));
    InMux I__1944 (
            .O(N__7903),
            .I(N__7878));
    InMux I__1943 (
            .O(N__7900),
            .I(N__7878));
    Span4Mux_h I__1942 (
            .O(N__7897),
            .I(N__7873));
    LocalMux I__1941 (
            .O(N__7892),
            .I(N__7873));
    InMux I__1940 (
            .O(N__7889),
            .I(N__7870));
    LocalMux I__1939 (
            .O(N__7886),
            .I(N__7867));
    InMux I__1938 (
            .O(N__7883),
            .I(N__7864));
    LocalMux I__1937 (
            .O(N__7878),
            .I(N__7857));
    Span4Mux_s2_v I__1936 (
            .O(N__7873),
            .I(N__7857));
    LocalMux I__1935 (
            .O(N__7870),
            .I(N__7857));
    Span4Mux_v I__1934 (
            .O(N__7867),
            .I(N__7854));
    LocalMux I__1933 (
            .O(N__7864),
            .I(N__7849));
    Span4Mux_v I__1932 (
            .O(N__7857),
            .I(N__7849));
    Odrv4 I__1931 (
            .O(N__7854),
            .I(acc_out_4));
    Odrv4 I__1930 (
            .O(N__7849),
            .I(acc_out_4));
    IoInMux I__1929 (
            .O(N__7844),
            .I(N__7841));
    LocalMux I__1928 (
            .O(N__7841),
            .I(N__7838));
    Odrv12 I__1927 (
            .O(N__7838),
            .I(out_c_4));
    InMux I__1926 (
            .O(N__7835),
            .I(N__7830));
    InMux I__1925 (
            .O(N__7834),
            .I(N__7825));
    InMux I__1924 (
            .O(N__7833),
            .I(N__7825));
    LocalMux I__1923 (
            .O(N__7830),
            .I(N__7822));
    LocalMux I__1922 (
            .O(N__7825),
            .I(N__7819));
    Span4Mux_h I__1921 (
            .O(N__7822),
            .I(N__7816));
    Odrv4 I__1920 (
            .O(N__7819),
            .I(b_reg_out_3));
    Odrv4 I__1919 (
            .O(N__7816),
            .I(b_reg_out_3));
    CEMux I__1918 (
            .O(N__7811),
            .I(N__7808));
    LocalMux I__1917 (
            .O(N__7808),
            .I(N__7805));
    Span4Mux_h I__1916 (
            .O(N__7805),
            .I(N__7800));
    CEMux I__1915 (
            .O(N__7804),
            .I(N__7797));
    CEMux I__1914 (
            .O(N__7803),
            .I(N__7794));
    Span4Mux_s2_v I__1913 (
            .O(N__7800),
            .I(N__7788));
    LocalMux I__1912 (
            .O(N__7797),
            .I(N__7788));
    LocalMux I__1911 (
            .O(N__7794),
            .I(N__7785));
    CEMux I__1910 (
            .O(N__7793),
            .I(N__7782));
    Span4Mux_v I__1909 (
            .O(N__7788),
            .I(N__7778));
    Span4Mux_v I__1908 (
            .O(N__7785),
            .I(N__7773));
    LocalMux I__1907 (
            .O(N__7782),
            .I(N__7773));
    CEMux I__1906 (
            .O(N__7781),
            .I(N__7770));
    Span4Mux_s2_v I__1905 (
            .O(N__7778),
            .I(N__7767));
    Span4Mux_h I__1904 (
            .O(N__7773),
            .I(N__7764));
    LocalMux I__1903 (
            .O(N__7770),
            .I(N__7761));
    Odrv4 I__1902 (
            .O(N__7767),
            .I(seq_B_LD_0_i));
    Odrv4 I__1901 (
            .O(N__7764),
            .I(seq_B_LD_0_i));
    Odrv4 I__1900 (
            .O(N__7761),
            .I(seq_B_LD_0_i));
    InMux I__1899 (
            .O(N__7754),
            .I(N__7751));
    LocalMux I__1898 (
            .O(N__7751),
            .I(N__7745));
    InMux I__1897 (
            .O(N__7750),
            .I(N__7742));
    InMux I__1896 (
            .O(N__7749),
            .I(N__7737));
    InMux I__1895 (
            .O(N__7748),
            .I(N__7734));
    Span4Mux_v I__1894 (
            .O(N__7745),
            .I(N__7729));
    LocalMux I__1893 (
            .O(N__7742),
            .I(N__7729));
    InMux I__1892 (
            .O(N__7741),
            .I(N__7726));
    InMux I__1891 (
            .O(N__7740),
            .I(N__7723));
    LocalMux I__1890 (
            .O(N__7737),
            .I(N__7720));
    LocalMux I__1889 (
            .O(N__7734),
            .I(N__7717));
    Span4Mux_v I__1888 (
            .O(N__7729),
            .I(N__7714));
    LocalMux I__1887 (
            .O(N__7726),
            .I(N__7711));
    LocalMux I__1886 (
            .O(N__7723),
            .I(N__7706));
    Span4Mux_s1_h I__1885 (
            .O(N__7720),
            .I(N__7706));
    Span12Mux_v I__1884 (
            .O(N__7717),
            .I(N__7703));
    Span4Mux_h I__1883 (
            .O(N__7714),
            .I(N__7700));
    Span4Mux_h I__1882 (
            .O(N__7711),
            .I(N__7697));
    Span4Mux_v I__1881 (
            .O(N__7706),
            .I(N__7694));
    Odrv12 I__1880 (
            .O(N__7703),
            .I(\pc.tbuf.g0_0_0 ));
    Odrv4 I__1879 (
            .O(N__7700),
            .I(\pc.tbuf.g0_0_0 ));
    Odrv4 I__1878 (
            .O(N__7697),
            .I(\pc.tbuf.g0_0_0 ));
    Odrv4 I__1877 (
            .O(N__7694),
            .I(\pc.tbuf.g0_0_0 ));
    InMux I__1876 (
            .O(N__7685),
            .I(N__7682));
    LocalMux I__1875 (
            .O(N__7682),
            .I(N__7675));
    InMux I__1874 (
            .O(N__7681),
            .I(N__7672));
    InMux I__1873 (
            .O(N__7680),
            .I(N__7669));
    InMux I__1872 (
            .O(N__7679),
            .I(N__7666));
    InMux I__1871 (
            .O(N__7678),
            .I(N__7663));
    Span4Mux_v I__1870 (
            .O(N__7675),
            .I(N__7660));
    LocalMux I__1869 (
            .O(N__7672),
            .I(N__7657));
    LocalMux I__1868 (
            .O(N__7669),
            .I(N__7654));
    LocalMux I__1867 (
            .O(N__7666),
            .I(N__7649));
    LocalMux I__1866 (
            .O(N__7663),
            .I(N__7649));
    Span4Mux_h I__1865 (
            .O(N__7660),
            .I(N__7646));
    Span4Mux_v I__1864 (
            .O(N__7657),
            .I(N__7643));
    Span4Mux_v I__1863 (
            .O(N__7654),
            .I(N__7638));
    Span4Mux_h I__1862 (
            .O(N__7649),
            .I(N__7638));
    Odrv4 I__1861 (
            .O(N__7646),
            .I(\pc.tbuf.g0Z0Z_3 ));
    Odrv4 I__1860 (
            .O(N__7643),
            .I(\pc.tbuf.g0Z0Z_3 ));
    Odrv4 I__1859 (
            .O(N__7638),
            .I(\pc.tbuf.g0Z0Z_3 ));
    CascadeMux I__1858 (
            .O(N__7631),
            .I(N__7627));
    CascadeMux I__1857 (
            .O(N__7630),
            .I(N__7624));
    InMux I__1856 (
            .O(N__7627),
            .I(N__7621));
    InMux I__1855 (
            .O(N__7624),
            .I(N__7615));
    LocalMux I__1854 (
            .O(N__7621),
            .I(N__7612));
    CascadeMux I__1853 (
            .O(N__7620),
            .I(N__7609));
    CascadeMux I__1852 (
            .O(N__7619),
            .I(N__7606));
    InMux I__1851 (
            .O(N__7618),
            .I(N__7603));
    LocalMux I__1850 (
            .O(N__7615),
            .I(N__7600));
    Span4Mux_v I__1849 (
            .O(N__7612),
            .I(N__7597));
    InMux I__1848 (
            .O(N__7609),
            .I(N__7594));
    InMux I__1847 (
            .O(N__7606),
            .I(N__7590));
    LocalMux I__1846 (
            .O(N__7603),
            .I(N__7587));
    Span4Mux_v I__1845 (
            .O(N__7600),
            .I(N__7584));
    Sp12to4 I__1844 (
            .O(N__7597),
            .I(N__7579));
    LocalMux I__1843 (
            .O(N__7594),
            .I(N__7579));
    CascadeMux I__1842 (
            .O(N__7593),
            .I(N__7576));
    LocalMux I__1841 (
            .O(N__7590),
            .I(N__7573));
    Span4Mux_v I__1840 (
            .O(N__7587),
            .I(N__7570));
    Span4Mux_h I__1839 (
            .O(N__7584),
            .I(N__7567));
    Span12Mux_s10_h I__1838 (
            .O(N__7579),
            .I(N__7564));
    InMux I__1837 (
            .O(N__7576),
            .I(N__7561));
    Span4Mux_v I__1836 (
            .O(N__7573),
            .I(N__7556));
    Span4Mux_v I__1835 (
            .O(N__7570),
            .I(N__7556));
    Odrv4 I__1834 (
            .O(N__7567),
            .I(\pc.tbuf.gZ0Z2 ));
    Odrv12 I__1833 (
            .O(N__7564),
            .I(\pc.tbuf.gZ0Z2 ));
    LocalMux I__1832 (
            .O(N__7561),
            .I(\pc.tbuf.gZ0Z2 ));
    Odrv4 I__1831 (
            .O(N__7556),
            .I(\pc.tbuf.gZ0Z2 ));
    InMux I__1830 (
            .O(N__7547),
            .I(N__7541));
    InMux I__1829 (
            .O(N__7546),
            .I(N__7537));
    InMux I__1828 (
            .O(N__7545),
            .I(N__7534));
    InMux I__1827 (
            .O(N__7544),
            .I(N__7531));
    LocalMux I__1826 (
            .O(N__7541),
            .I(N__7528));
    InMux I__1825 (
            .O(N__7540),
            .I(N__7525));
    LocalMux I__1824 (
            .O(N__7537),
            .I(N__7521));
    LocalMux I__1823 (
            .O(N__7534),
            .I(N__7518));
    LocalMux I__1822 (
            .O(N__7531),
            .I(N__7515));
    Span4Mux_v I__1821 (
            .O(N__7528),
            .I(N__7510));
    LocalMux I__1820 (
            .O(N__7525),
            .I(N__7510));
    InMux I__1819 (
            .O(N__7524),
            .I(N__7507));
    Span4Mux_h I__1818 (
            .O(N__7521),
            .I(N__7500));
    Span4Mux_s3_h I__1817 (
            .O(N__7518),
            .I(N__7500));
    Span4Mux_s3_h I__1816 (
            .O(N__7515),
            .I(N__7500));
    Odrv4 I__1815 (
            .O(N__7510),
            .I(alu_out_m_1_3));
    LocalMux I__1814 (
            .O(N__7507),
            .I(alu_out_m_1_3));
    Odrv4 I__1813 (
            .O(N__7500),
            .I(alu_out_m_1_3));
    IoInMux I__1812 (
            .O(N__7493),
            .I(N__7490));
    LocalMux I__1811 (
            .O(N__7490),
            .I(N__7487));
    Odrv12 I__1810 (
            .O(N__7487),
            .I(out_c_3));
    CEMux I__1809 (
            .O(N__7484),
            .I(N__7481));
    LocalMux I__1808 (
            .O(N__7481),
            .I(N__7470));
    CEMux I__1807 (
            .O(N__7480),
            .I(N__7467));
    InMux I__1806 (
            .O(N__7479),
            .I(N__7464));
    CEMux I__1805 (
            .O(N__7478),
            .I(N__7461));
    InMux I__1804 (
            .O(N__7477),
            .I(N__7458));
    InMux I__1803 (
            .O(N__7476),
            .I(N__7451));
    CEMux I__1802 (
            .O(N__7475),
            .I(N__7448));
    CEMux I__1801 (
            .O(N__7474),
            .I(N__7445));
    CEMux I__1800 (
            .O(N__7473),
            .I(N__7442));
    Span4Mux_v I__1799 (
            .O(N__7470),
            .I(N__7438));
    LocalMux I__1798 (
            .O(N__7467),
            .I(N__7435));
    LocalMux I__1797 (
            .O(N__7464),
            .I(N__7432));
    LocalMux I__1796 (
            .O(N__7461),
            .I(N__7427));
    LocalMux I__1795 (
            .O(N__7458),
            .I(N__7427));
    InMux I__1794 (
            .O(N__7457),
            .I(N__7424));
    InMux I__1793 (
            .O(N__7456),
            .I(N__7419));
    InMux I__1792 (
            .O(N__7455),
            .I(N__7419));
    InMux I__1791 (
            .O(N__7454),
            .I(N__7416));
    LocalMux I__1790 (
            .O(N__7451),
            .I(N__7413));
    LocalMux I__1789 (
            .O(N__7448),
            .I(N__7409));
    LocalMux I__1788 (
            .O(N__7445),
            .I(N__7404));
    LocalMux I__1787 (
            .O(N__7442),
            .I(N__7404));
    InMux I__1786 (
            .O(N__7441),
            .I(N__7401));
    Span4Mux_h I__1785 (
            .O(N__7438),
            .I(N__7389));
    Span4Mux_v I__1784 (
            .O(N__7435),
            .I(N__7389));
    Span4Mux_v I__1783 (
            .O(N__7432),
            .I(N__7389));
    Span4Mux_h I__1782 (
            .O(N__7427),
            .I(N__7389));
    LocalMux I__1781 (
            .O(N__7424),
            .I(N__7385));
    LocalMux I__1780 (
            .O(N__7419),
            .I(N__7378));
    LocalMux I__1779 (
            .O(N__7416),
            .I(N__7378));
    Span4Mux_v I__1778 (
            .O(N__7413),
            .I(N__7378));
    InMux I__1777 (
            .O(N__7412),
            .I(N__7375));
    Span4Mux_h I__1776 (
            .O(N__7409),
            .I(N__7370));
    Span4Mux_v I__1775 (
            .O(N__7404),
            .I(N__7370));
    LocalMux I__1774 (
            .O(N__7401),
            .I(N__7367));
    InMux I__1773 (
            .O(N__7400),
            .I(N__7364));
    InMux I__1772 (
            .O(N__7399),
            .I(N__7361));
    InMux I__1771 (
            .O(N__7398),
            .I(N__7358));
    Span4Mux_h I__1770 (
            .O(N__7389),
            .I(N__7355));
    InMux I__1769 (
            .O(N__7388),
            .I(N__7352));
    Span4Mux_s2_v I__1768 (
            .O(N__7385),
            .I(N__7345));
    Span4Mux_v I__1767 (
            .O(N__7378),
            .I(N__7345));
    LocalMux I__1766 (
            .O(N__7375),
            .I(N__7345));
    Span4Mux_h I__1765 (
            .O(N__7370),
            .I(N__7340));
    Span4Mux_v I__1764 (
            .O(N__7367),
            .I(N__7340));
    LocalMux I__1763 (
            .O(N__7364),
            .I(N__7333));
    LocalMux I__1762 (
            .O(N__7361),
            .I(N__7333));
    LocalMux I__1761 (
            .O(N__7358),
            .I(N__7333));
    Odrv4 I__1760 (
            .O(N__7355),
            .I(OUT_LD));
    LocalMux I__1759 (
            .O(N__7352),
            .I(OUT_LD));
    Odrv4 I__1758 (
            .O(N__7345),
            .I(OUT_LD));
    Odrv4 I__1757 (
            .O(N__7340),
            .I(OUT_LD));
    Odrv12 I__1756 (
            .O(N__7333),
            .I(OUT_LD));
    SRMux I__1755 (
            .O(N__7322),
            .I(N__7214));
    SRMux I__1754 (
            .O(N__7321),
            .I(N__7214));
    SRMux I__1753 (
            .O(N__7320),
            .I(N__7214));
    SRMux I__1752 (
            .O(N__7319),
            .I(N__7214));
    SRMux I__1751 (
            .O(N__7318),
            .I(N__7214));
    SRMux I__1750 (
            .O(N__7317),
            .I(N__7214));
    SRMux I__1749 (
            .O(N__7316),
            .I(N__7214));
    SRMux I__1748 (
            .O(N__7315),
            .I(N__7214));
    SRMux I__1747 (
            .O(N__7314),
            .I(N__7214));
    SRMux I__1746 (
            .O(N__7313),
            .I(N__7214));
    SRMux I__1745 (
            .O(N__7312),
            .I(N__7214));
    SRMux I__1744 (
            .O(N__7311),
            .I(N__7214));
    SRMux I__1743 (
            .O(N__7310),
            .I(N__7214));
    SRMux I__1742 (
            .O(N__7309),
            .I(N__7214));
    SRMux I__1741 (
            .O(N__7308),
            .I(N__7214));
    SRMux I__1740 (
            .O(N__7307),
            .I(N__7214));
    SRMux I__1739 (
            .O(N__7306),
            .I(N__7214));
    SRMux I__1738 (
            .O(N__7305),
            .I(N__7214));
    SRMux I__1737 (
            .O(N__7304),
            .I(N__7214));
    SRMux I__1736 (
            .O(N__7303),
            .I(N__7214));
    SRMux I__1735 (
            .O(N__7302),
            .I(N__7214));
    SRMux I__1734 (
            .O(N__7301),
            .I(N__7214));
    SRMux I__1733 (
            .O(N__7300),
            .I(N__7214));
    SRMux I__1732 (
            .O(N__7299),
            .I(N__7214));
    SRMux I__1731 (
            .O(N__7298),
            .I(N__7214));
    SRMux I__1730 (
            .O(N__7297),
            .I(N__7214));
    SRMux I__1729 (
            .O(N__7296),
            .I(N__7214));
    SRMux I__1728 (
            .O(N__7295),
            .I(N__7214));
    SRMux I__1727 (
            .O(N__7294),
            .I(N__7214));
    SRMux I__1726 (
            .O(N__7293),
            .I(N__7214));
    SRMux I__1725 (
            .O(N__7292),
            .I(N__7214));
    SRMux I__1724 (
            .O(N__7291),
            .I(N__7214));
    SRMux I__1723 (
            .O(N__7290),
            .I(N__7214));
    SRMux I__1722 (
            .O(N__7289),
            .I(N__7214));
    SRMux I__1721 (
            .O(N__7288),
            .I(N__7214));
    SRMux I__1720 (
            .O(N__7287),
            .I(N__7214));
    GlobalMux I__1719 (
            .O(N__7214),
            .I(N__7211));
    gio2CtrlBuf I__1718 (
            .O(N__7211),
            .I(clr_c_g));
    CascadeMux I__1717 (
            .O(N__7208),
            .I(mem_data_2_7_0__N_29_mux_cascade_));
    IoInMux I__1716 (
            .O(N__7205),
            .I(N__7202));
    LocalMux I__1715 (
            .O(N__7202),
            .I(N__7199));
    Odrv12 I__1714 (
            .O(N__7199),
            .I(out_c_6));
    CascadeMux I__1713 (
            .O(N__7196),
            .I(N__7193));
    InMux I__1712 (
            .O(N__7193),
            .I(N__7187));
    InMux I__1711 (
            .O(N__7192),
            .I(N__7187));
    LocalMux I__1710 (
            .O(N__7187),
            .I(N__7183));
    InMux I__1709 (
            .O(N__7186),
            .I(N__7180));
    Span4Mux_v I__1708 (
            .O(N__7183),
            .I(N__7168));
    LocalMux I__1707 (
            .O(N__7180),
            .I(N__7168));
    InMux I__1706 (
            .O(N__7179),
            .I(N__7156));
    InMux I__1705 (
            .O(N__7178),
            .I(N__7156));
    InMux I__1704 (
            .O(N__7177),
            .I(N__7156));
    InMux I__1703 (
            .O(N__7176),
            .I(N__7156));
    InMux I__1702 (
            .O(N__7175),
            .I(N__7156));
    InMux I__1701 (
            .O(N__7174),
            .I(N__7151));
    InMux I__1700 (
            .O(N__7173),
            .I(N__7151));
    Span4Mux_h I__1699 (
            .O(N__7168),
            .I(N__7148));
    InMux I__1698 (
            .O(N__7167),
            .I(N__7145));
    LocalMux I__1697 (
            .O(N__7156),
            .I(N__7142));
    LocalMux I__1696 (
            .O(N__7151),
            .I(N__7139));
    Odrv4 I__1695 (
            .O(N__7148),
            .I(mar_out_2));
    LocalMux I__1694 (
            .O(N__7145),
            .I(mar_out_2));
    Odrv4 I__1693 (
            .O(N__7142),
            .I(mar_out_2));
    Odrv12 I__1692 (
            .O(N__7139),
            .I(mar_out_2));
    InMux I__1691 (
            .O(N__7130),
            .I(N__7122));
    InMux I__1690 (
            .O(N__7129),
            .I(N__7122));
    CascadeMux I__1689 (
            .O(N__7128),
            .I(N__7115));
    CascadeMux I__1688 (
            .O(N__7127),
            .I(N__7110));
    LocalMux I__1687 (
            .O(N__7122),
            .I(N__7105));
    InMux I__1686 (
            .O(N__7121),
            .I(N__7102));
    InMux I__1685 (
            .O(N__7120),
            .I(N__7099));
    InMux I__1684 (
            .O(N__7119),
            .I(N__7094));
    InMux I__1683 (
            .O(N__7118),
            .I(N__7094));
    InMux I__1682 (
            .O(N__7115),
            .I(N__7083));
    InMux I__1681 (
            .O(N__7114),
            .I(N__7083));
    InMux I__1680 (
            .O(N__7113),
            .I(N__7083));
    InMux I__1679 (
            .O(N__7110),
            .I(N__7083));
    InMux I__1678 (
            .O(N__7109),
            .I(N__7083));
    InMux I__1677 (
            .O(N__7108),
            .I(N__7080));
    Span4Mux_v I__1676 (
            .O(N__7105),
            .I(N__7077));
    LocalMux I__1675 (
            .O(N__7102),
            .I(N__7070));
    LocalMux I__1674 (
            .O(N__7099),
            .I(N__7070));
    LocalMux I__1673 (
            .O(N__7094),
            .I(N__7070));
    LocalMux I__1672 (
            .O(N__7083),
            .I(N__7067));
    LocalMux I__1671 (
            .O(N__7080),
            .I(mar_out_1));
    Odrv4 I__1670 (
            .O(N__7077),
            .I(mar_out_1));
    Odrv12 I__1669 (
            .O(N__7070),
            .I(mar_out_1));
    Odrv4 I__1668 (
            .O(N__7067),
            .I(mar_out_1));
    CascadeMux I__1667 (
            .O(N__7058),
            .I(N__7054));
    InMux I__1666 (
            .O(N__7057),
            .I(N__7048));
    InMux I__1665 (
            .O(N__7054),
            .I(N__7048));
    CascadeMux I__1664 (
            .O(N__7053),
            .I(N__7039));
    LocalMux I__1663 (
            .O(N__7048),
            .I(N__7036));
    CascadeMux I__1662 (
            .O(N__7047),
            .I(N__7033));
    CascadeMux I__1661 (
            .O(N__7046),
            .I(N__7030));
    CascadeMux I__1660 (
            .O(N__7045),
            .I(N__7025));
    InMux I__1659 (
            .O(N__7044),
            .I(N__7022));
    CascadeMux I__1658 (
            .O(N__7043),
            .I(N__7019));
    CascadeMux I__1657 (
            .O(N__7042),
            .I(N__7015));
    InMux I__1656 (
            .O(N__7039),
            .I(N__7012));
    Span4Mux_h I__1655 (
            .O(N__7036),
            .I(N__7009));
    InMux I__1654 (
            .O(N__7033),
            .I(N__6998));
    InMux I__1653 (
            .O(N__7030),
            .I(N__6998));
    InMux I__1652 (
            .O(N__7029),
            .I(N__6998));
    InMux I__1651 (
            .O(N__7028),
            .I(N__6998));
    InMux I__1650 (
            .O(N__7025),
            .I(N__6998));
    LocalMux I__1649 (
            .O(N__7022),
            .I(N__6995));
    InMux I__1648 (
            .O(N__7019),
            .I(N__6988));
    InMux I__1647 (
            .O(N__7018),
            .I(N__6988));
    InMux I__1646 (
            .O(N__7015),
            .I(N__6988));
    LocalMux I__1645 (
            .O(N__7012),
            .I(N__6985));
    Span4Mux_h I__1644 (
            .O(N__7009),
            .I(N__6980));
    LocalMux I__1643 (
            .O(N__6998),
            .I(N__6980));
    Span12Mux_s10_v I__1642 (
            .O(N__6995),
            .I(N__6975));
    LocalMux I__1641 (
            .O(N__6988),
            .I(N__6975));
    Odrv4 I__1640 (
            .O(N__6985),
            .I(mar_out_3));
    Odrv4 I__1639 (
            .O(N__6980),
            .I(mar_out_3));
    Odrv12 I__1638 (
            .O(N__6975),
            .I(mar_out_3));
    InMux I__1637 (
            .O(N__6968),
            .I(N__6957));
    InMux I__1636 (
            .O(N__6967),
            .I(N__6952));
    InMux I__1635 (
            .O(N__6966),
            .I(N__6952));
    InMux I__1634 (
            .O(N__6965),
            .I(N__6949));
    InMux I__1633 (
            .O(N__6964),
            .I(N__6938));
    InMux I__1632 (
            .O(N__6963),
            .I(N__6938));
    InMux I__1631 (
            .O(N__6962),
            .I(N__6938));
    InMux I__1630 (
            .O(N__6961),
            .I(N__6938));
    InMux I__1629 (
            .O(N__6960),
            .I(N__6938));
    LocalMux I__1628 (
            .O(N__6957),
            .I(N__6935));
    LocalMux I__1627 (
            .O(N__6952),
            .I(N__6927));
    LocalMux I__1626 (
            .O(N__6949),
            .I(N__6927));
    LocalMux I__1625 (
            .O(N__6938),
            .I(N__6924));
    Span4Mux_v I__1624 (
            .O(N__6935),
            .I(N__6921));
    InMux I__1623 (
            .O(N__6934),
            .I(N__6914));
    InMux I__1622 (
            .O(N__6933),
            .I(N__6914));
    InMux I__1621 (
            .O(N__6932),
            .I(N__6914));
    Span4Mux_v I__1620 (
            .O(N__6927),
            .I(N__6909));
    Span4Mux_h I__1619 (
            .O(N__6924),
            .I(N__6909));
    Odrv4 I__1618 (
            .O(N__6921),
            .I(mar_out_0));
    LocalMux I__1617 (
            .O(N__6914),
            .I(mar_out_0));
    Odrv4 I__1616 (
            .O(N__6909),
            .I(mar_out_0));
    InMux I__1615 (
            .O(N__6902),
            .I(N__6895));
    InMux I__1614 (
            .O(N__6901),
            .I(N__6895));
    InMux I__1613 (
            .O(N__6900),
            .I(N__6892));
    LocalMux I__1612 (
            .O(N__6895),
            .I(N__6887));
    LocalMux I__1611 (
            .O(N__6892),
            .I(N__6884));
    CascadeMux I__1610 (
            .O(N__6891),
            .I(N__6881));
    CascadeMux I__1609 (
            .O(N__6890),
            .I(N__6878));
    Span4Mux_s2_h I__1608 (
            .O(N__6887),
            .I(N__6875));
    Span4Mux_h I__1607 (
            .O(N__6884),
            .I(N__6872));
    InMux I__1606 (
            .O(N__6881),
            .I(N__6869));
    InMux I__1605 (
            .O(N__6878),
            .I(N__6866));
    Span4Mux_h I__1604 (
            .O(N__6875),
            .I(N__6863));
    Odrv4 I__1603 (
            .O(N__6872),
            .I(mem_data_2_7_0__i2_mux_0));
    LocalMux I__1602 (
            .O(N__6869),
            .I(mem_data_2_7_0__i2_mux_0));
    LocalMux I__1601 (
            .O(N__6866),
            .I(mem_data_2_7_0__i2_mux_0));
    Odrv4 I__1600 (
            .O(N__6863),
            .I(mem_data_2_7_0__i2_mux_0));
    InMux I__1599 (
            .O(N__6854),
            .I(N__6851));
    LocalMux I__1598 (
            .O(N__6851),
            .I(N__6848));
    Span4Mux_h I__1597 (
            .O(N__6848),
            .I(N__6844));
    InMux I__1596 (
            .O(N__6847),
            .I(N__6841));
    Odrv4 I__1595 (
            .O(N__6844),
            .I(b_reg_out_1));
    LocalMux I__1594 (
            .O(N__6841),
            .I(b_reg_out_1));
    CascadeMux I__1593 (
            .O(N__6836),
            .I(N__6833));
    InMux I__1592 (
            .O(N__6833),
            .I(N__6830));
    LocalMux I__1591 (
            .O(N__6830),
            .I(N__6826));
    InMux I__1590 (
            .O(N__6829),
            .I(N__6823));
    Span4Mux_s3_v I__1589 (
            .O(N__6826),
            .I(N__6817));
    LocalMux I__1588 (
            .O(N__6823),
            .I(N__6814));
    InMux I__1587 (
            .O(N__6822),
            .I(N__6811));
    InMux I__1586 (
            .O(N__6821),
            .I(N__6808));
    InMux I__1585 (
            .O(N__6820),
            .I(N__6805));
    Span4Mux_s1_h I__1584 (
            .O(N__6817),
            .I(N__6800));
    Span4Mux_s3_v I__1583 (
            .O(N__6814),
            .I(N__6800));
    LocalMux I__1582 (
            .O(N__6811),
            .I(acc_out_m_6));
    LocalMux I__1581 (
            .O(N__6808),
            .I(acc_out_m_6));
    LocalMux I__1580 (
            .O(N__6805),
            .I(acc_out_m_6));
    Odrv4 I__1579 (
            .O(N__6800),
            .I(acc_out_m_6));
    InMux I__1578 (
            .O(N__6791),
            .I(N__6786));
    InMux I__1577 (
            .O(N__6790),
            .I(N__6783));
    InMux I__1576 (
            .O(N__6789),
            .I(N__6779));
    LocalMux I__1575 (
            .O(N__6786),
            .I(N__6775));
    LocalMux I__1574 (
            .O(N__6783),
            .I(N__6772));
    InMux I__1573 (
            .O(N__6782),
            .I(N__6769));
    LocalMux I__1572 (
            .O(N__6779),
            .I(N__6766));
    InMux I__1571 (
            .O(N__6778),
            .I(N__6763));
    Span4Mux_s3_v I__1570 (
            .O(N__6775),
            .I(N__6756));
    Span4Mux_s3_v I__1569 (
            .O(N__6772),
            .I(N__6756));
    LocalMux I__1568 (
            .O(N__6769),
            .I(N__6756));
    Span4Mux_s3_h I__1567 (
            .O(N__6766),
            .I(N__6753));
    LocalMux I__1566 (
            .O(N__6763),
            .I(alu_out_m_6));
    Odrv4 I__1565 (
            .O(N__6756),
            .I(alu_out_m_6));
    Odrv4 I__1564 (
            .O(N__6753),
            .I(alu_out_m_6));
    CascadeMux I__1563 (
            .O(N__6746),
            .I(N__6742));
    InMux I__1562 (
            .O(N__6745),
            .I(N__6739));
    InMux I__1561 (
            .O(N__6742),
            .I(N__6736));
    LocalMux I__1560 (
            .O(N__6739),
            .I(N__6729));
    LocalMux I__1559 (
            .O(N__6736),
            .I(N__6729));
    CascadeMux I__1558 (
            .O(N__6735),
            .I(N__6726));
    CascadeMux I__1557 (
            .O(N__6734),
            .I(N__6723));
    Span4Mux_v I__1556 (
            .O(N__6729),
            .I(N__6720));
    InMux I__1555 (
            .O(N__6726),
            .I(N__6717));
    InMux I__1554 (
            .O(N__6723),
            .I(N__6714));
    Span4Mux_h I__1553 (
            .O(N__6720),
            .I(N__6711));
    LocalMux I__1552 (
            .O(N__6717),
            .I(mem_data_2_7_0__N_29_mux));
    LocalMux I__1551 (
            .O(N__6714),
            .I(mem_data_2_7_0__N_29_mux));
    Odrv4 I__1550 (
            .O(N__6711),
            .I(mem_data_2_7_0__N_29_mux));
    InMux I__1549 (
            .O(N__6704),
            .I(N__6700));
    InMux I__1548 (
            .O(N__6703),
            .I(N__6697));
    LocalMux I__1547 (
            .O(N__6700),
            .I(b_reg_out_6));
    LocalMux I__1546 (
            .O(N__6697),
            .I(b_reg_out_6));
    InMux I__1545 (
            .O(N__6692),
            .I(N__6687));
    InMux I__1544 (
            .O(N__6691),
            .I(N__6684));
    CascadeMux I__1543 (
            .O(N__6690),
            .I(N__6680));
    LocalMux I__1542 (
            .O(N__6687),
            .I(N__6677));
    LocalMux I__1541 (
            .O(N__6684),
            .I(N__6674));
    InMux I__1540 (
            .O(N__6683),
            .I(N__6671));
    InMux I__1539 (
            .O(N__6680),
            .I(N__6667));
    Span4Mux_v I__1538 (
            .O(N__6677),
            .I(N__6664));
    Span4Mux_s2_v I__1537 (
            .O(N__6674),
            .I(N__6661));
    LocalMux I__1536 (
            .O(N__6671),
            .I(N__6658));
    InMux I__1535 (
            .O(N__6670),
            .I(N__6655));
    LocalMux I__1534 (
            .O(N__6667),
            .I(N__6652));
    Odrv4 I__1533 (
            .O(N__6664),
            .I(acc_out_m_5));
    Odrv4 I__1532 (
            .O(N__6661),
            .I(acc_out_m_5));
    Odrv4 I__1531 (
            .O(N__6658),
            .I(acc_out_m_5));
    LocalMux I__1530 (
            .O(N__6655),
            .I(acc_out_m_5));
    Odrv12 I__1529 (
            .O(N__6652),
            .I(acc_out_m_5));
    InMux I__1528 (
            .O(N__6641),
            .I(N__6638));
    LocalMux I__1527 (
            .O(N__6638),
            .I(N__6631));
    InMux I__1526 (
            .O(N__6637),
            .I(N__6628));
    InMux I__1525 (
            .O(N__6636),
            .I(N__6625));
    InMux I__1524 (
            .O(N__6635),
            .I(N__6622));
    InMux I__1523 (
            .O(N__6634),
            .I(N__6619));
    Span4Mux_h I__1522 (
            .O(N__6631),
            .I(N__6610));
    LocalMux I__1521 (
            .O(N__6628),
            .I(N__6610));
    LocalMux I__1520 (
            .O(N__6625),
            .I(N__6610));
    LocalMux I__1519 (
            .O(N__6622),
            .I(N__6610));
    LocalMux I__1518 (
            .O(N__6619),
            .I(alu_out_m_5));
    Odrv4 I__1517 (
            .O(N__6610),
            .I(alu_out_m_5));
    CascadeMux I__1516 (
            .O(N__6605),
            .I(N__6601));
    CascadeMux I__1515 (
            .O(N__6604),
            .I(N__6595));
    InMux I__1514 (
            .O(N__6601),
            .I(N__6592));
    InMux I__1513 (
            .O(N__6600),
            .I(N__6589));
    CascadeMux I__1512 (
            .O(N__6599),
            .I(N__6586));
    CascadeMux I__1511 (
            .O(N__6598),
            .I(N__6583));
    InMux I__1510 (
            .O(N__6595),
            .I(N__6580));
    LocalMux I__1509 (
            .O(N__6592),
            .I(N__6575));
    LocalMux I__1508 (
            .O(N__6589),
            .I(N__6575));
    InMux I__1507 (
            .O(N__6586),
            .I(N__6572));
    InMux I__1506 (
            .O(N__6583),
            .I(N__6569));
    LocalMux I__1505 (
            .O(N__6580),
            .I(N__6564));
    Span4Mux_h I__1504 (
            .O(N__6575),
            .I(N__6564));
    LocalMux I__1503 (
            .O(N__6572),
            .I(m20));
    LocalMux I__1502 (
            .O(N__6569),
            .I(m20));
    Odrv4 I__1501 (
            .O(N__6564),
            .I(m20));
    InMux I__1500 (
            .O(N__6557),
            .I(N__6548));
    InMux I__1499 (
            .O(N__6556),
            .I(N__6543));
    InMux I__1498 (
            .O(N__6555),
            .I(N__6543));
    InMux I__1497 (
            .O(N__6554),
            .I(N__6538));
    InMux I__1496 (
            .O(N__6553),
            .I(N__6538));
    InMux I__1495 (
            .O(N__6552),
            .I(N__6531));
    InMux I__1494 (
            .O(N__6551),
            .I(N__6528));
    LocalMux I__1493 (
            .O(N__6548),
            .I(N__6514));
    LocalMux I__1492 (
            .O(N__6543),
            .I(N__6514));
    LocalMux I__1491 (
            .O(N__6538),
            .I(N__6514));
    InMux I__1490 (
            .O(N__6537),
            .I(N__6511));
    InMux I__1489 (
            .O(N__6536),
            .I(N__6504));
    InMux I__1488 (
            .O(N__6535),
            .I(N__6504));
    InMux I__1487 (
            .O(N__6534),
            .I(N__6504));
    LocalMux I__1486 (
            .O(N__6531),
            .I(N__6499));
    LocalMux I__1485 (
            .O(N__6528),
            .I(N__6499));
    InMux I__1484 (
            .O(N__6527),
            .I(N__6496));
    InMux I__1483 (
            .O(N__6526),
            .I(N__6489));
    InMux I__1482 (
            .O(N__6525),
            .I(N__6489));
    InMux I__1481 (
            .O(N__6524),
            .I(N__6489));
    InMux I__1480 (
            .O(N__6523),
            .I(N__6486));
    InMux I__1479 (
            .O(N__6522),
            .I(N__6483));
    InMux I__1478 (
            .O(N__6521),
            .I(N__6479));
    Span4Mux_v I__1477 (
            .O(N__6514),
            .I(N__6474));
    LocalMux I__1476 (
            .O(N__6511),
            .I(N__6474));
    LocalMux I__1475 (
            .O(N__6504),
            .I(N__6467));
    Span4Mux_s2_v I__1474 (
            .O(N__6499),
            .I(N__6467));
    LocalMux I__1473 (
            .O(N__6496),
            .I(N__6467));
    LocalMux I__1472 (
            .O(N__6489),
            .I(N__6460));
    LocalMux I__1471 (
            .O(N__6486),
            .I(N__6455));
    LocalMux I__1470 (
            .O(N__6483),
            .I(N__6455));
    InMux I__1469 (
            .O(N__6482),
            .I(N__6452));
    LocalMux I__1468 (
            .O(N__6479),
            .I(N__6445));
    Span4Mux_h I__1467 (
            .O(N__6474),
            .I(N__6445));
    Span4Mux_h I__1466 (
            .O(N__6467),
            .I(N__6445));
    InMux I__1465 (
            .O(N__6466),
            .I(N__6438));
    InMux I__1464 (
            .O(N__6465),
            .I(N__6438));
    InMux I__1463 (
            .O(N__6464),
            .I(N__6438));
    InMux I__1462 (
            .O(N__6463),
            .I(N__6435));
    Odrv12 I__1461 (
            .O(N__6460),
            .I(ROM_OE));
    Odrv4 I__1460 (
            .O(N__6455),
            .I(ROM_OE));
    LocalMux I__1459 (
            .O(N__6452),
            .I(ROM_OE));
    Odrv4 I__1458 (
            .O(N__6445),
            .I(ROM_OE));
    LocalMux I__1457 (
            .O(N__6438),
            .I(ROM_OE));
    LocalMux I__1456 (
            .O(N__6435),
            .I(ROM_OE));
    IoInMux I__1455 (
            .O(N__6422),
            .I(N__6419));
    LocalMux I__1454 (
            .O(N__6419),
            .I(N__6416));
    Span4Mux_s1_v I__1453 (
            .O(N__6416),
            .I(N__6413));
    Span4Mux_h I__1452 (
            .O(N__6413),
            .I(N__6410));
    Odrv4 I__1451 (
            .O(N__6410),
            .I(out_c_5));
    IoInMux I__1450 (
            .O(N__6407),
            .I(N__6404));
    LocalMux I__1449 (
            .O(N__6404),
            .I(N__6401));
    Odrv12 I__1448 (
            .O(N__6401),
            .I(out_c_2));
    IoInMux I__1447 (
            .O(N__6398),
            .I(N__6395));
    LocalMux I__1446 (
            .O(N__6395),
            .I(N__6392));
    IoSpan4Mux I__1445 (
            .O(N__6392),
            .I(N__6389));
    Span4Mux_s1_h I__1444 (
            .O(N__6389),
            .I(N__6386));
    Odrv4 I__1443 (
            .O(N__6386),
            .I(out_c_0));
    CEMux I__1442 (
            .O(N__6383),
            .I(N__6379));
    CEMux I__1441 (
            .O(N__6382),
            .I(N__6376));
    LocalMux I__1440 (
            .O(N__6379),
            .I(N__6373));
    LocalMux I__1439 (
            .O(N__6376),
            .I(N__6370));
    Span4Mux_v I__1438 (
            .O(N__6373),
            .I(N__6365));
    Span4Mux_v I__1437 (
            .O(N__6370),
            .I(N__6365));
    Span4Mux_h I__1436 (
            .O(N__6365),
            .I(N__6362));
    Odrv4 I__1435 (
            .O(N__6362),
            .I(\mar.MAR_LD_0_0 ));
    InMux I__1434 (
            .O(N__6359),
            .I(N__6353));
    InMux I__1433 (
            .O(N__6358),
            .I(N__6353));
    LocalMux I__1432 (
            .O(N__6353),
            .I(b_reg_out_5));
    InMux I__1431 (
            .O(N__6350),
            .I(N__6347));
    LocalMux I__1430 (
            .O(N__6347),
            .I(N__6343));
    InMux I__1429 (
            .O(N__6346),
            .I(N__6340));
    Span4Mux_h I__1428 (
            .O(N__6343),
            .I(N__6335));
    LocalMux I__1427 (
            .O(N__6340),
            .I(N__6335));
    Span4Mux_v I__1426 (
            .O(N__6335),
            .I(N__6331));
    InMux I__1425 (
            .O(N__6334),
            .I(N__6328));
    Span4Mux_h I__1424 (
            .O(N__6331),
            .I(N__6324));
    LocalMux I__1423 (
            .O(N__6328),
            .I(N__6321));
    InMux I__1422 (
            .O(N__6327),
            .I(N__6318));
    Odrv4 I__1421 (
            .O(N__6324),
            .I(acc_out_m_7));
    Odrv12 I__1420 (
            .O(N__6321),
            .I(acc_out_m_7));
    LocalMux I__1419 (
            .O(N__6318),
            .I(acc_out_m_7));
    InMux I__1418 (
            .O(N__6311),
            .I(N__6306));
    InMux I__1417 (
            .O(N__6310),
            .I(N__6303));
    CascadeMux I__1416 (
            .O(N__6309),
            .I(N__6300));
    LocalMux I__1415 (
            .O(N__6306),
            .I(N__6297));
    LocalMux I__1414 (
            .O(N__6303),
            .I(N__6294));
    InMux I__1413 (
            .O(N__6300),
            .I(N__6290));
    Span4Mux_h I__1412 (
            .O(N__6297),
            .I(N__6285));
    Span4Mux_v I__1411 (
            .O(N__6294),
            .I(N__6285));
    InMux I__1410 (
            .O(N__6293),
            .I(N__6282));
    LocalMux I__1409 (
            .O(N__6290),
            .I(N__6279));
    Span4Mux_h I__1408 (
            .O(N__6285),
            .I(N__6276));
    LocalMux I__1407 (
            .O(N__6282),
            .I(alu_out_m_7));
    Odrv12 I__1406 (
            .O(N__6279),
            .I(alu_out_m_7));
    Odrv4 I__1405 (
            .O(N__6276),
            .I(alu_out_m_7));
    InMux I__1404 (
            .O(N__6269),
            .I(N__6265));
    CascadeMux I__1403 (
            .O(N__6268),
            .I(N__6262));
    LocalMux I__1402 (
            .O(N__6265),
            .I(N__6259));
    InMux I__1401 (
            .O(N__6262),
            .I(N__6256));
    Span4Mux_v I__1400 (
            .O(N__6259),
            .I(N__6251));
    LocalMux I__1399 (
            .O(N__6256),
            .I(N__6251));
    Span4Mux_h I__1398 (
            .O(N__6251),
            .I(N__6248));
    Odrv4 I__1397 (
            .O(N__6248),
            .I(b_reg_out_7));
    InMux I__1396 (
            .O(N__6245),
            .I(N__6240));
    InMux I__1395 (
            .O(N__6244),
            .I(N__6235));
    InMux I__1394 (
            .O(N__6243),
            .I(N__6235));
    LocalMux I__1393 (
            .O(N__6240),
            .I(N__6232));
    LocalMux I__1392 (
            .O(N__6235),
            .I(N__6229));
    Odrv12 I__1391 (
            .O(N__6232),
            .I(b_reg_out_0));
    Odrv4 I__1390 (
            .O(N__6229),
            .I(b_reg_out_0));
    CascadeMux I__1389 (
            .O(N__6224),
            .I(\mem.i2_mux_cascade_ ));
    InMux I__1388 (
            .O(N__6221),
            .I(N__6218));
    LocalMux I__1387 (
            .O(N__6218),
            .I(N__6215));
    Span4Mux_h I__1386 (
            .O(N__6215),
            .I(N__6212));
    Odrv4 I__1385 (
            .O(N__6212),
            .I(\pc.N_7 ));
    InMux I__1384 (
            .O(N__6209),
            .I(N__6206));
    LocalMux I__1383 (
            .O(N__6206),
            .I(N__6202));
    InMux I__1382 (
            .O(N__6205),
            .I(N__6199));
    Odrv4 I__1381 (
            .O(N__6202),
            .I(b_reg_out_4));
    LocalMux I__1380 (
            .O(N__6199),
            .I(b_reg_out_4));
    InMux I__1379 (
            .O(N__6194),
            .I(N__6187));
    InMux I__1378 (
            .O(N__6193),
            .I(N__6183));
    InMux I__1377 (
            .O(N__6192),
            .I(N__6180));
    InMux I__1376 (
            .O(N__6191),
            .I(N__6175));
    InMux I__1375 (
            .O(N__6190),
            .I(N__6175));
    LocalMux I__1374 (
            .O(N__6187),
            .I(N__6172));
    InMux I__1373 (
            .O(N__6186),
            .I(N__6169));
    LocalMux I__1372 (
            .O(N__6183),
            .I(N__6153));
    LocalMux I__1371 (
            .O(N__6180),
            .I(N__6148));
    LocalMux I__1370 (
            .O(N__6175),
            .I(N__6148));
    Span4Mux_v I__1369 (
            .O(N__6172),
            .I(N__6143));
    LocalMux I__1368 (
            .O(N__6169),
            .I(N__6143));
    InMux I__1367 (
            .O(N__6168),
            .I(N__6136));
    InMux I__1366 (
            .O(N__6167),
            .I(N__6136));
    InMux I__1365 (
            .O(N__6166),
            .I(N__6136));
    InMux I__1364 (
            .O(N__6165),
            .I(N__6131));
    InMux I__1363 (
            .O(N__6164),
            .I(N__6131));
    InMux I__1362 (
            .O(N__6163),
            .I(N__6124));
    InMux I__1361 (
            .O(N__6162),
            .I(N__6124));
    InMux I__1360 (
            .O(N__6161),
            .I(N__6124));
    InMux I__1359 (
            .O(N__6160),
            .I(N__6119));
    InMux I__1358 (
            .O(N__6159),
            .I(N__6119));
    InMux I__1357 (
            .O(N__6158),
            .I(N__6112));
    InMux I__1356 (
            .O(N__6157),
            .I(N__6112));
    InMux I__1355 (
            .O(N__6156),
            .I(N__6112));
    Odrv12 I__1354 (
            .O(N__6153),
            .I(seq_S0_0));
    Odrv4 I__1353 (
            .O(N__6148),
            .I(seq_S0_0));
    Odrv4 I__1352 (
            .O(N__6143),
            .I(seq_S0_0));
    LocalMux I__1351 (
            .O(N__6136),
            .I(seq_S0_0));
    LocalMux I__1350 (
            .O(N__6131),
            .I(seq_S0_0));
    LocalMux I__1349 (
            .O(N__6124),
            .I(seq_S0_0));
    LocalMux I__1348 (
            .O(N__6119),
            .I(seq_S0_0));
    LocalMux I__1347 (
            .O(N__6112),
            .I(seq_S0_0));
    CascadeMux I__1346 (
            .O(N__6095),
            .I(N__6092));
    InMux I__1345 (
            .O(N__6092),
            .I(N__6089));
    LocalMux I__1344 (
            .O(N__6089),
            .I(\ALU_main.N_45 ));
    InMux I__1343 (
            .O(N__6086),
            .I(N__6083));
    LocalMux I__1342 (
            .O(N__6083),
            .I(N__6080));
    Span4Mux_h I__1341 (
            .O(N__6080),
            .I(N__6076));
    InMux I__1340 (
            .O(N__6079),
            .I(N__6073));
    Odrv4 I__1339 (
            .O(N__6076),
            .I(bus_5));
    LocalMux I__1338 (
            .O(N__6073),
            .I(bus_5));
    InMux I__1337 (
            .O(N__6068),
            .I(N__6064));
    InMux I__1336 (
            .O(N__6067),
            .I(N__6061));
    LocalMux I__1335 (
            .O(N__6064),
            .I(N__6055));
    LocalMux I__1334 (
            .O(N__6061),
            .I(N__6055));
    InMux I__1333 (
            .O(N__6060),
            .I(N__6052));
    Span4Mux_v I__1332 (
            .O(N__6055),
            .I(N__6045));
    LocalMux I__1331 (
            .O(N__6052),
            .I(N__6045));
    InMux I__1330 (
            .O(N__6051),
            .I(N__6042));
    InMux I__1329 (
            .O(N__6050),
            .I(N__6039));
    Span4Mux_h I__1328 (
            .O(N__6045),
            .I(N__6036));
    LocalMux I__1327 (
            .O(N__6042),
            .I(acc_out_0));
    LocalMux I__1326 (
            .O(N__6039),
            .I(acc_out_0));
    Odrv4 I__1325 (
            .O(N__6036),
            .I(acc_out_0));
    InMux I__1324 (
            .O(N__6029),
            .I(N__6025));
    InMux I__1323 (
            .O(N__6028),
            .I(N__6021));
    LocalMux I__1322 (
            .O(N__6025),
            .I(N__6018));
    InMux I__1321 (
            .O(N__6024),
            .I(N__6015));
    LocalMux I__1320 (
            .O(N__6021),
            .I(N__6011));
    Span4Mux_v I__1319 (
            .O(N__6018),
            .I(N__6006));
    LocalMux I__1318 (
            .O(N__6015),
            .I(N__6006));
    InMux I__1317 (
            .O(N__6014),
            .I(N__6003));
    Span4Mux_h I__1316 (
            .O(N__6011),
            .I(N__6000));
    Odrv4 I__1315 (
            .O(N__6006),
            .I(acc_out_1));
    LocalMux I__1314 (
            .O(N__6003),
            .I(acc_out_1));
    Odrv4 I__1313 (
            .O(N__6000),
            .I(acc_out_1));
    CascadeMux I__1312 (
            .O(N__5993),
            .I(N__5986));
    InMux I__1311 (
            .O(N__5992),
            .I(N__5979));
    InMux I__1310 (
            .O(N__5991),
            .I(N__5979));
    InMux I__1309 (
            .O(N__5990),
            .I(N__5979));
    InMux I__1308 (
            .O(N__5989),
            .I(N__5976));
    InMux I__1307 (
            .O(N__5986),
            .I(N__5973));
    LocalMux I__1306 (
            .O(N__5979),
            .I(N__5970));
    LocalMux I__1305 (
            .O(N__5976),
            .I(N__5967));
    LocalMux I__1304 (
            .O(N__5973),
            .I(N__5964));
    Span4Mux_h I__1303 (
            .O(N__5970),
            .I(N__5961));
    Span4Mux_v I__1302 (
            .O(N__5967),
            .I(N__5958));
    Span4Mux_v I__1301 (
            .O(N__5964),
            .I(N__5955));
    Odrv4 I__1300 (
            .O(N__5961),
            .I(acc_out_2));
    Odrv4 I__1299 (
            .O(N__5958),
            .I(acc_out_2));
    Odrv4 I__1298 (
            .O(N__5955),
            .I(acc_out_2));
    CEMux I__1297 (
            .O(N__5948),
            .I(N__5944));
    CEMux I__1296 (
            .O(N__5947),
            .I(N__5941));
    LocalMux I__1295 (
            .O(N__5944),
            .I(N__5938));
    LocalMux I__1294 (
            .O(N__5941),
            .I(N__5935));
    Span4Mux_v I__1293 (
            .O(N__5938),
            .I(N__5932));
    Span4Mux_h I__1292 (
            .O(N__5935),
            .I(N__5929));
    Odrv4 I__1291 (
            .O(N__5932),
            .I(seq_ACC_LD_0_i));
    Odrv4 I__1290 (
            .O(N__5929),
            .I(seq_ACC_LD_0_i));
    CascadeMux I__1289 (
            .O(N__5924),
            .I(N__5921));
    InMux I__1288 (
            .O(N__5921),
            .I(N__5918));
    LocalMux I__1287 (
            .O(N__5918),
            .I(N__5915));
    Odrv4 I__1286 (
            .O(N__5915),
            .I(\ALU_main.N_47 ));
    CascadeMux I__1285 (
            .O(N__5912),
            .I(N__5909));
    InMux I__1284 (
            .O(N__5909),
            .I(N__5903));
    InMux I__1283 (
            .O(N__5908),
            .I(N__5900));
    InMux I__1282 (
            .O(N__5907),
            .I(N__5895));
    InMux I__1281 (
            .O(N__5906),
            .I(N__5895));
    LocalMux I__1280 (
            .O(N__5903),
            .I(N__5892));
    LocalMux I__1279 (
            .O(N__5900),
            .I(acc_out_6));
    LocalMux I__1278 (
            .O(N__5895),
            .I(acc_out_6));
    Odrv4 I__1277 (
            .O(N__5892),
            .I(acc_out_6));
    InMux I__1276 (
            .O(N__5885),
            .I(N__5882));
    LocalMux I__1275 (
            .O(N__5882),
            .I(N__5879));
    Odrv4 I__1274 (
            .O(N__5879),
            .I(\ALU_main.un1_A_axb_6_l_ofxZ0 ));
    InMux I__1273 (
            .O(N__5876),
            .I(N__5870));
    InMux I__1272 (
            .O(N__5875),
            .I(N__5870));
    LocalMux I__1271 (
            .O(N__5870),
            .I(N__5867));
    Span4Mux_h I__1270 (
            .O(N__5867),
            .I(N__5863));
    InMux I__1269 (
            .O(N__5866),
            .I(N__5860));
    Odrv4 I__1268 (
            .O(N__5863),
            .I(acc_out_7));
    LocalMux I__1267 (
            .O(N__5860),
            .I(acc_out_7));
    CascadeMux I__1266 (
            .O(N__5855),
            .I(N__5849));
    InMux I__1265 (
            .O(N__5854),
            .I(N__5842));
    InMux I__1264 (
            .O(N__5853),
            .I(N__5842));
    InMux I__1263 (
            .O(N__5852),
            .I(N__5842));
    InMux I__1262 (
            .O(N__5849),
            .I(N__5839));
    LocalMux I__1261 (
            .O(N__5842),
            .I(N__5834));
    LocalMux I__1260 (
            .O(N__5839),
            .I(N__5834));
    Span4Mux_h I__1259 (
            .O(N__5834),
            .I(N__5831));
    Odrv4 I__1258 (
            .O(N__5831),
            .I(acc_out_5));
    CascadeMux I__1257 (
            .O(N__5828),
            .I(N__5824));
    InMux I__1256 (
            .O(N__5827),
            .I(N__5817));
    InMux I__1255 (
            .O(N__5824),
            .I(N__5814));
    InMux I__1254 (
            .O(N__5823),
            .I(N__5811));
    InMux I__1253 (
            .O(N__5822),
            .I(N__5808));
    InMux I__1252 (
            .O(N__5821),
            .I(N__5803));
    InMux I__1251 (
            .O(N__5820),
            .I(N__5803));
    LocalMux I__1250 (
            .O(N__5817),
            .I(N__5800));
    LocalMux I__1249 (
            .O(N__5814),
            .I(N__5797));
    LocalMux I__1248 (
            .O(N__5811),
            .I(N__5794));
    LocalMux I__1247 (
            .O(N__5808),
            .I(N__5789));
    LocalMux I__1246 (
            .O(N__5803),
            .I(N__5789));
    Span4Mux_h I__1245 (
            .O(N__5800),
            .I(N__5784));
    Span4Mux_h I__1244 (
            .O(N__5797),
            .I(N__5784));
    Odrv4 I__1243 (
            .O(N__5794),
            .I(acc_out_3));
    Odrv4 I__1242 (
            .O(N__5789),
            .I(acc_out_3));
    Odrv4 I__1241 (
            .O(N__5784),
            .I(acc_out_3));
    InMux I__1240 (
            .O(N__5777),
            .I(N__5774));
    LocalMux I__1239 (
            .O(N__5774),
            .I(N__5771));
    Odrv4 I__1238 (
            .O(N__5771),
            .I(\ALU_main.un1_A_cry_3_c_RNI552PZ0Z2 ));
    InMux I__1237 (
            .O(N__5768),
            .I(N__5764));
    InMux I__1236 (
            .O(N__5767),
            .I(N__5757));
    LocalMux I__1235 (
            .O(N__5764),
            .I(N__5754));
    InMux I__1234 (
            .O(N__5763),
            .I(N__5749));
    InMux I__1233 (
            .O(N__5762),
            .I(N__5749));
    InMux I__1232 (
            .O(N__5761),
            .I(N__5743));
    InMux I__1231 (
            .O(N__5760),
            .I(N__5738));
    LocalMux I__1230 (
            .O(N__5757),
            .I(N__5735));
    Span4Mux_v I__1229 (
            .O(N__5754),
            .I(N__5732));
    LocalMux I__1228 (
            .O(N__5749),
            .I(N__5729));
    InMux I__1227 (
            .O(N__5748),
            .I(N__5722));
    InMux I__1226 (
            .O(N__5747),
            .I(N__5722));
    InMux I__1225 (
            .O(N__5746),
            .I(N__5722));
    LocalMux I__1224 (
            .O(N__5743),
            .I(N__5719));
    InMux I__1223 (
            .O(N__5742),
            .I(N__5714));
    InMux I__1222 (
            .O(N__5741),
            .I(N__5714));
    LocalMux I__1221 (
            .O(N__5738),
            .I(N__5711));
    Span4Mux_s3_v I__1220 (
            .O(N__5735),
            .I(N__5702));
    Span4Mux_h I__1219 (
            .O(N__5732),
            .I(N__5702));
    Span4Mux_v I__1218 (
            .O(N__5729),
            .I(N__5702));
    LocalMux I__1217 (
            .O(N__5722),
            .I(N__5702));
    Span4Mux_h I__1216 (
            .O(N__5719),
            .I(N__5697));
    LocalMux I__1215 (
            .O(N__5714),
            .I(N__5697));
    Span12Mux_s10_h I__1214 (
            .O(N__5711),
            .I(N__5694));
    Span4Mux_h I__1213 (
            .O(N__5702),
            .I(N__5689));
    Span4Mux_v I__1212 (
            .O(N__5697),
            .I(N__5689));
    Odrv12 I__1211 (
            .O(N__5694),
            .I(seq_un1_ALU_en_0));
    Odrv4 I__1210 (
            .O(N__5689),
            .I(seq_un1_ALU_en_0));
    CascadeMux I__1209 (
            .O(N__5684),
            .I(N__5676));
    InMux I__1208 (
            .O(N__5683),
            .I(N__5668));
    InMux I__1207 (
            .O(N__5682),
            .I(N__5668));
    InMux I__1206 (
            .O(N__5681),
            .I(N__5665));
    InMux I__1205 (
            .O(N__5680),
            .I(N__5662));
    InMux I__1204 (
            .O(N__5679),
            .I(N__5659));
    InMux I__1203 (
            .O(N__5676),
            .I(N__5656));
    InMux I__1202 (
            .O(N__5675),
            .I(N__5653));
    InMux I__1201 (
            .O(N__5674),
            .I(N__5648));
    InMux I__1200 (
            .O(N__5673),
            .I(N__5648));
    LocalMux I__1199 (
            .O(N__5668),
            .I(N__5645));
    LocalMux I__1198 (
            .O(N__5665),
            .I(N__5640));
    LocalMux I__1197 (
            .O(N__5662),
            .I(N__5637));
    LocalMux I__1196 (
            .O(N__5659),
            .I(N__5634));
    LocalMux I__1195 (
            .O(N__5656),
            .I(N__5631));
    LocalMux I__1194 (
            .O(N__5653),
            .I(N__5626));
    LocalMux I__1193 (
            .O(N__5648),
            .I(N__5626));
    Span4Mux_v I__1192 (
            .O(N__5645),
            .I(N__5623));
    InMux I__1191 (
            .O(N__5644),
            .I(N__5618));
    InMux I__1190 (
            .O(N__5643),
            .I(N__5618));
    Span4Mux_v I__1189 (
            .O(N__5640),
            .I(N__5611));
    Span4Mux_h I__1188 (
            .O(N__5637),
            .I(N__5611));
    Span4Mux_v I__1187 (
            .O(N__5634),
            .I(N__5611));
    Span4Mux_h I__1186 (
            .O(N__5631),
            .I(N__5602));
    Span4Mux_h I__1185 (
            .O(N__5626),
            .I(N__5602));
    Span4Mux_h I__1184 (
            .O(N__5623),
            .I(N__5602));
    LocalMux I__1183 (
            .O(N__5618),
            .I(N__5602));
    Odrv4 I__1182 (
            .O(N__5611),
            .I(seq_S1_0));
    Odrv4 I__1181 (
            .O(N__5602),
            .I(seq_S1_0));
    CascadeMux I__1180 (
            .O(N__5597),
            .I(alu_out_m_4_cascade_));
    InMux I__1179 (
            .O(N__5594),
            .I(N__5591));
    LocalMux I__1178 (
            .O(N__5591),
            .I(N__5587));
    InMux I__1177 (
            .O(N__5590),
            .I(N__5584));
    Span4Mux_s1_h I__1176 (
            .O(N__5587),
            .I(N__5581));
    LocalMux I__1175 (
            .O(N__5584),
            .I(N__5578));
    Span4Mux_h I__1174 (
            .O(N__5581),
            .I(N__5575));
    Span4Mux_v I__1173 (
            .O(N__5578),
            .I(N__5572));
    Odrv4 I__1172 (
            .O(N__5575),
            .I(bus_4));
    Odrv4 I__1171 (
            .O(N__5572),
            .I(bus_4));
    CascadeMux I__1170 (
            .O(N__5567),
            .I(bus_4_cascade_));
    InMux I__1169 (
            .O(N__5564),
            .I(N__5558));
    InMux I__1168 (
            .O(N__5563),
            .I(N__5555));
    InMux I__1167 (
            .O(N__5562),
            .I(N__5550));
    InMux I__1166 (
            .O(N__5561),
            .I(N__5550));
    LocalMux I__1165 (
            .O(N__5558),
            .I(N__5542));
    LocalMux I__1164 (
            .O(N__5555),
            .I(N__5539));
    LocalMux I__1163 (
            .O(N__5550),
            .I(N__5536));
    InMux I__1162 (
            .O(N__5549),
            .I(N__5531));
    InMux I__1161 (
            .O(N__5548),
            .I(N__5531));
    InMux I__1160 (
            .O(N__5547),
            .I(N__5526));
    InMux I__1159 (
            .O(N__5546),
            .I(N__5526));
    InMux I__1158 (
            .O(N__5545),
            .I(N__5523));
    Odrv4 I__1157 (
            .O(N__5542),
            .I(ir_out_4));
    Odrv12 I__1156 (
            .O(N__5539),
            .I(ir_out_4));
    Odrv4 I__1155 (
            .O(N__5536),
            .I(ir_out_4));
    LocalMux I__1154 (
            .O(N__5531),
            .I(ir_out_4));
    LocalMux I__1153 (
            .O(N__5526),
            .I(ir_out_4));
    LocalMux I__1152 (
            .O(N__5523),
            .I(ir_out_4));
    InMux I__1151 (
            .O(N__5510),
            .I(N__5507));
    LocalMux I__1150 (
            .O(N__5507),
            .I(N_4_0));
    InMux I__1149 (
            .O(N__5504),
            .I(N__5501));
    LocalMux I__1148 (
            .O(N__5501),
            .I(N__5491));
    InMux I__1147 (
            .O(N__5500),
            .I(N__5488));
    InMux I__1146 (
            .O(N__5499),
            .I(N__5483));
    InMux I__1145 (
            .O(N__5498),
            .I(N__5483));
    InMux I__1144 (
            .O(N__5497),
            .I(N__5478));
    InMux I__1143 (
            .O(N__5496),
            .I(N__5478));
    InMux I__1142 (
            .O(N__5495),
            .I(N__5475));
    InMux I__1141 (
            .O(N__5494),
            .I(N__5472));
    Span4Mux_v I__1140 (
            .O(N__5491),
            .I(N__5469));
    LocalMux I__1139 (
            .O(N__5488),
            .I(ir_out_i_2_5));
    LocalMux I__1138 (
            .O(N__5483),
            .I(ir_out_i_2_5));
    LocalMux I__1137 (
            .O(N__5478),
            .I(ir_out_i_2_5));
    LocalMux I__1136 (
            .O(N__5475),
            .I(ir_out_i_2_5));
    LocalMux I__1135 (
            .O(N__5472),
            .I(ir_out_i_2_5));
    Odrv4 I__1134 (
            .O(N__5469),
            .I(ir_out_i_2_5));
    InMux I__1133 (
            .O(N__5456),
            .I(N__5452));
    InMux I__1132 (
            .O(N__5455),
            .I(N__5449));
    LocalMux I__1131 (
            .O(N__5452),
            .I(N__5440));
    LocalMux I__1130 (
            .O(N__5449),
            .I(N__5437));
    InMux I__1129 (
            .O(N__5448),
            .I(N__5430));
    InMux I__1128 (
            .O(N__5447),
            .I(N__5430));
    InMux I__1127 (
            .O(N__5446),
            .I(N__5430));
    InMux I__1126 (
            .O(N__5445),
            .I(N__5427));
    InMux I__1125 (
            .O(N__5444),
            .I(N__5422));
    InMux I__1124 (
            .O(N__5443),
            .I(N__5422));
    Span4Mux_h I__1123 (
            .O(N__5440),
            .I(N__5419));
    Odrv12 I__1122 (
            .O(N__5437),
            .I(ir_out_4_rep1));
    LocalMux I__1121 (
            .O(N__5430),
            .I(ir_out_4_rep1));
    LocalMux I__1120 (
            .O(N__5427),
            .I(ir_out_4_rep1));
    LocalMux I__1119 (
            .O(N__5422),
            .I(ir_out_4_rep1));
    Odrv4 I__1118 (
            .O(N__5419),
            .I(ir_out_4_rep1));
    InMux I__1117 (
            .O(N__5408),
            .I(N__5402));
    CascadeMux I__1116 (
            .O(N__5407),
            .I(N__5399));
    InMux I__1115 (
            .O(N__5406),
            .I(N__5394));
    InMux I__1114 (
            .O(N__5405),
            .I(N__5391));
    LocalMux I__1113 (
            .O(N__5402),
            .I(N__5388));
    InMux I__1112 (
            .O(N__5399),
            .I(N__5385));
    InMux I__1111 (
            .O(N__5398),
            .I(N__5380));
    InMux I__1110 (
            .O(N__5397),
            .I(N__5380));
    LocalMux I__1109 (
            .O(N__5394),
            .I(N__5377));
    LocalMux I__1108 (
            .O(N__5391),
            .I(IR_ff7_q_0_fast));
    Odrv4 I__1107 (
            .O(N__5388),
            .I(IR_ff7_q_0_fast));
    LocalMux I__1106 (
            .O(N__5385),
            .I(IR_ff7_q_0_fast));
    LocalMux I__1105 (
            .O(N__5380),
            .I(IR_ff7_q_0_fast));
    Odrv4 I__1104 (
            .O(N__5377),
            .I(IR_ff7_q_0_fast));
    InMux I__1103 (
            .O(N__5366),
            .I(N__5359));
    InMux I__1102 (
            .O(N__5365),
            .I(N__5354));
    InMux I__1101 (
            .O(N__5364),
            .I(N__5354));
    InMux I__1100 (
            .O(N__5363),
            .I(N__5351));
    CascadeMux I__1099 (
            .O(N__5362),
            .I(N__5347));
    LocalMux I__1098 (
            .O(N__5359),
            .I(N__5342));
    LocalMux I__1097 (
            .O(N__5354),
            .I(N__5342));
    LocalMux I__1096 (
            .O(N__5351),
            .I(N__5339));
    InMux I__1095 (
            .O(N__5350),
            .I(N__5334));
    InMux I__1094 (
            .O(N__5347),
            .I(N__5334));
    Span4Mux_v I__1093 (
            .O(N__5342),
            .I(N__5327));
    Span4Mux_h I__1092 (
            .O(N__5339),
            .I(N__5327));
    LocalMux I__1091 (
            .O(N__5334),
            .I(N__5327));
    Span4Mux_h I__1090 (
            .O(N__5327),
            .I(N__5322));
    InMux I__1089 (
            .O(N__5326),
            .I(N__5317));
    InMux I__1088 (
            .O(N__5325),
            .I(N__5317));
    Odrv4 I__1087 (
            .O(N__5322),
            .I(\seq.counter.TZ0Z_4 ));
    LocalMux I__1086 (
            .O(N__5317),
            .I(\seq.counter.TZ0Z_4 ));
    InMux I__1085 (
            .O(N__5312),
            .I(N__5306));
    InMux I__1084 (
            .O(N__5311),
            .I(N__5303));
    InMux I__1083 (
            .O(N__5310),
            .I(N__5300));
    InMux I__1082 (
            .O(N__5309),
            .I(N__5296));
    LocalMux I__1081 (
            .O(N__5306),
            .I(N__5292));
    LocalMux I__1080 (
            .O(N__5303),
            .I(N__5285));
    LocalMux I__1079 (
            .O(N__5300),
            .I(N__5285));
    CascadeMux I__1078 (
            .O(N__5299),
            .I(N__5282));
    LocalMux I__1077 (
            .O(N__5296),
            .I(N__5278));
    InMux I__1076 (
            .O(N__5295),
            .I(N__5275));
    Span4Mux_h I__1075 (
            .O(N__5292),
            .I(N__5272));
    InMux I__1074 (
            .O(N__5291),
            .I(N__5267));
    InMux I__1073 (
            .O(N__5290),
            .I(N__5267));
    Span4Mux_h I__1072 (
            .O(N__5285),
            .I(N__5264));
    InMux I__1071 (
            .O(N__5282),
            .I(N__5259));
    InMux I__1070 (
            .O(N__5281),
            .I(N__5259));
    Odrv4 I__1069 (
            .O(N__5278),
            .I(ir_out_7));
    LocalMux I__1068 (
            .O(N__5275),
            .I(ir_out_7));
    Odrv4 I__1067 (
            .O(N__5272),
            .I(ir_out_7));
    LocalMux I__1066 (
            .O(N__5267),
            .I(ir_out_7));
    Odrv4 I__1065 (
            .O(N__5264),
            .I(ir_out_7));
    LocalMux I__1064 (
            .O(N__5259),
            .I(ir_out_7));
    CascadeMux I__1063 (
            .O(N__5246),
            .I(\seq.g0_i_a3_0Z0Z_2_cascade_ ));
    InMux I__1062 (
            .O(N__5243),
            .I(N__5240));
    LocalMux I__1061 (
            .O(N__5240),
            .I(N__5237));
    Span4Mux_h I__1060 (
            .O(N__5237),
            .I(N__5234));
    Odrv4 I__1059 (
            .O(N__5234),
            .I(\seq.g0_i_a3Z0Z_2 ));
    CascadeMux I__1058 (
            .O(N__5231),
            .I(seq_S0_0_cascade_));
    InMux I__1057 (
            .O(N__5228),
            .I(N__5225));
    LocalMux I__1056 (
            .O(N__5225),
            .I(\ALU_main.un1_A_axb_5_l_ofxZ0 ));
    InMux I__1055 (
            .O(N__5222),
            .I(N__5219));
    LocalMux I__1054 (
            .O(N__5219),
            .I(N__5213));
    InMux I__1053 (
            .O(N__5218),
            .I(N__5210));
    InMux I__1052 (
            .O(N__5217),
            .I(N__5207));
    InMux I__1051 (
            .O(N__5216),
            .I(N__5204));
    Span4Mux_s3_v I__1050 (
            .O(N__5213),
            .I(N__5197));
    LocalMux I__1049 (
            .O(N__5210),
            .I(N__5197));
    LocalMux I__1048 (
            .O(N__5207),
            .I(N__5192));
    LocalMux I__1047 (
            .O(N__5204),
            .I(N__5192));
    InMux I__1046 (
            .O(N__5203),
            .I(N__5189));
    CascadeMux I__1045 (
            .O(N__5202),
            .I(N__5185));
    Span4Mux_v I__1044 (
            .O(N__5197),
            .I(N__5182));
    Span4Mux_v I__1043 (
            .O(N__5192),
            .I(N__5179));
    LocalMux I__1042 (
            .O(N__5189),
            .I(N__5176));
    InMux I__1041 (
            .O(N__5188),
            .I(N__5173));
    InMux I__1040 (
            .O(N__5185),
            .I(N__5170));
    Span4Mux_s1_h I__1039 (
            .O(N__5182),
            .I(N__5165));
    Span4Mux_s1_h I__1038 (
            .O(N__5179),
            .I(N__5165));
    Odrv12 I__1037 (
            .O(N__5176),
            .I(\seq.counter.TZ0Z_3 ));
    LocalMux I__1036 (
            .O(N__5173),
            .I(\seq.counter.TZ0Z_3 ));
    LocalMux I__1035 (
            .O(N__5170),
            .I(\seq.counter.TZ0Z_3 ));
    Odrv4 I__1034 (
            .O(N__5165),
            .I(\seq.counter.TZ0Z_3 ));
    InMux I__1033 (
            .O(N__5156),
            .I(N__5151));
    InMux I__1032 (
            .O(N__5155),
            .I(N__5148));
    InMux I__1031 (
            .O(N__5154),
            .I(N__5144));
    LocalMux I__1030 (
            .O(N__5151),
            .I(N__5139));
    LocalMux I__1029 (
            .O(N__5148),
            .I(N__5139));
    CascadeMux I__1028 (
            .O(N__5147),
            .I(N__5135));
    LocalMux I__1027 (
            .O(N__5144),
            .I(N__5130));
    Span4Mux_h I__1026 (
            .O(N__5139),
            .I(N__5127));
    InMux I__1025 (
            .O(N__5138),
            .I(N__5120));
    InMux I__1024 (
            .O(N__5135),
            .I(N__5120));
    InMux I__1023 (
            .O(N__5134),
            .I(N__5120));
    InMux I__1022 (
            .O(N__5133),
            .I(N__5117));
    Odrv12 I__1021 (
            .O(N__5130),
            .I(\seq.D_2 ));
    Odrv4 I__1020 (
            .O(N__5127),
            .I(\seq.D_2 ));
    LocalMux I__1019 (
            .O(N__5120),
            .I(\seq.D_2 ));
    LocalMux I__1018 (
            .O(N__5117),
            .I(\seq.D_2 ));
    CascadeMux I__1017 (
            .O(N__5108),
            .I(N__5105));
    InMux I__1016 (
            .O(N__5105),
            .I(N__5102));
    LocalMux I__1015 (
            .O(N__5102),
            .I(N__5099));
    Odrv4 I__1014 (
            .O(N__5099),
            .I(\seq.B_LD_0_2_tz ));
    InMux I__1013 (
            .O(N__5096),
            .I(N__5093));
    LocalMux I__1012 (
            .O(N__5093),
            .I(N__5089));
    InMux I__1011 (
            .O(N__5092),
            .I(N__5085));
    Span4Mux_v I__1010 (
            .O(N__5089),
            .I(N__5082));
    InMux I__1009 (
            .O(N__5088),
            .I(N__5079));
    LocalMux I__1008 (
            .O(N__5085),
            .I(N__5075));
    Span4Mux_h I__1007 (
            .O(N__5082),
            .I(N__5070));
    LocalMux I__1006 (
            .O(N__5079),
            .I(N__5070));
    InMux I__1005 (
            .O(N__5078),
            .I(N__5067));
    Odrv12 I__1004 (
            .O(N__5075),
            .I(\seq.D_1 ));
    Odrv4 I__1003 (
            .O(N__5070),
            .I(\seq.D_1 ));
    LocalMux I__1002 (
            .O(N__5067),
            .I(\seq.D_1 ));
    CascadeMux I__1001 (
            .O(N__5060),
            .I(N__5057));
    InMux I__1000 (
            .O(N__5057),
            .I(N__5054));
    LocalMux I__999 (
            .O(N__5054),
            .I(\ALU_main.un1_A_axb_1_l_ofxZ0 ));
    InMux I__998 (
            .O(N__5051),
            .I(N__5048));
    LocalMux I__997 (
            .O(N__5048),
            .I(\ALU_main.un1_A_axb_4_l_ofxZ0 ));
    CascadeMux I__996 (
            .O(N__5045),
            .I(ALU_main_N_42_0_cascade_));
    InMux I__995 (
            .O(N__5042),
            .I(N__5039));
    LocalMux I__994 (
            .O(N__5039),
            .I(un1_A_cry_0_c_RNIPCLO2));
    CascadeMux I__993 (
            .O(N__5036),
            .I(ALU_main_N_41_0_cascade_));
    InMux I__992 (
            .O(N__5033),
            .I(N__5030));
    LocalMux I__991 (
            .O(N__5030),
            .I(N__5026));
    InMux I__990 (
            .O(N__5029),
            .I(N__5023));
    Span4Mux_s3_h I__989 (
            .O(N__5026),
            .I(N__5020));
    LocalMux I__988 (
            .O(N__5023),
            .I(un1_A_cry_0_s));
    Odrv4 I__987 (
            .O(N__5020),
            .I(un1_A_cry_0_s));
    InMux I__986 (
            .O(N__5015),
            .I(N__5009));
    InMux I__985 (
            .O(N__5014),
            .I(N__5009));
    LocalMux I__984 (
            .O(N__5009),
            .I(N__5006));
    Span4Mux_h I__983 (
            .O(N__5006),
            .I(N__4999));
    InMux I__982 (
            .O(N__5005),
            .I(N__4992));
    InMux I__981 (
            .O(N__5004),
            .I(N__4992));
    InMux I__980 (
            .O(N__5003),
            .I(N__4992));
    InMux I__979 (
            .O(N__5002),
            .I(N__4989));
    Odrv4 I__978 (
            .O(N__4999),
            .I(\seq.D_4 ));
    LocalMux I__977 (
            .O(N__4992),
            .I(\seq.D_4 ));
    LocalMux I__976 (
            .O(N__4989),
            .I(\seq.D_4 ));
    InMux I__975 (
            .O(N__4982),
            .I(N__4977));
    InMux I__974 (
            .O(N__4981),
            .I(N__4972));
    InMux I__973 (
            .O(N__4980),
            .I(N__4972));
    LocalMux I__972 (
            .O(N__4977),
            .I(N__4969));
    LocalMux I__971 (
            .O(N__4972),
            .I(N__4966));
    Span4Mux_v I__970 (
            .O(N__4969),
            .I(N__4958));
    Span4Mux_v I__969 (
            .O(N__4966),
            .I(N__4958));
    InMux I__968 (
            .O(N__4965),
            .I(N__4953));
    InMux I__967 (
            .O(N__4964),
            .I(N__4953));
    InMux I__966 (
            .O(N__4963),
            .I(N__4950));
    Odrv4 I__965 (
            .O(N__4958),
            .I(\seq.DZ0Z_0 ));
    LocalMux I__964 (
            .O(N__4953),
            .I(\seq.DZ0Z_0 ));
    LocalMux I__963 (
            .O(N__4950),
            .I(\seq.DZ0Z_0 ));
    CascadeMux I__962 (
            .O(N__4943),
            .I(N__4940));
    InMux I__961 (
            .O(N__4940),
            .I(N__4937));
    LocalMux I__960 (
            .O(N__4937),
            .I(N__4934));
    Span4Mux_h I__959 (
            .O(N__4934),
            .I(N__4931));
    Odrv4 I__958 (
            .O(N__4931),
            .I(\seq.g2Z0Z_1 ));
    CascadeMux I__957 (
            .O(N__4928),
            .I(N__4925));
    InMux I__956 (
            .O(N__4925),
            .I(N__4922));
    LocalMux I__955 (
            .O(N__4922),
            .I(\ALU_main.un1_A_axb_0_l_ofxZ0 ));
    InMux I__954 (
            .O(N__4919),
            .I(N__4916));
    LocalMux I__953 (
            .O(N__4916),
            .I(\ALU_main.un1_A_axb_3_l_ofxZ0 ));
    InMux I__952 (
            .O(N__4913),
            .I(N__4910));
    LocalMux I__951 (
            .O(N__4910),
            .I(\ALU_main.un1_A_cry_4_c_RNI9D6PZ0Z2 ));
    CascadeMux I__950 (
            .O(N__4907),
            .I(\ALU_main.N_46_cascade_ ));
    InMux I__949 (
            .O(N__4904),
            .I(N__4901));
    LocalMux I__948 (
            .O(N__4901),
            .I(N__4898));
    Span4Mux_v I__947 (
            .O(N__4898),
            .I(N__4894));
    InMux I__946 (
            .O(N__4897),
            .I(N__4891));
    Span4Mux_h I__945 (
            .O(N__4894),
            .I(N__4884));
    LocalMux I__944 (
            .O(N__4891),
            .I(N__4884));
    InMux I__943 (
            .O(N__4890),
            .I(N__4879));
    InMux I__942 (
            .O(N__4889),
            .I(N__4879));
    Odrv4 I__941 (
            .O(N__4884),
            .I(\seq.D_3 ));
    LocalMux I__940 (
            .O(N__4879),
            .I(\seq.D_3 ));
    CascadeMux I__939 (
            .O(N__4874),
            .I(\seq.counter.ACC_LD_0_0_cascade_ ));
    InMux I__938 (
            .O(N__4871),
            .I(N__4868));
    LocalMux I__937 (
            .O(N__4868),
            .I(N__4865));
    Odrv12 I__936 (
            .O(N__4865),
            .I(\pc.program_counter_m_0_1 ));
    InMux I__935 (
            .O(N__4862),
            .I(N__4859));
    LocalMux I__934 (
            .O(N__4859),
            .I(\pc.tbuf.out_1_1_ivZ0Z_0 ));
    CascadeMux I__933 (
            .O(N__4856),
            .I(mem_data_2_7_0__N_11_0_cascade_));
    InMux I__932 (
            .O(N__4853),
            .I(N__4850));
    LocalMux I__931 (
            .O(N__4850),
            .I(\pc.program_counter_4_rn_2_1 ));
    InMux I__930 (
            .O(N__4847),
            .I(N__4844));
    LocalMux I__929 (
            .O(N__4844),
            .I(\pc.program_counter_4_sn_1 ));
    CascadeMux I__928 (
            .O(N__4841),
            .I(\pc.g0_1_0_cascade_ ));
    CascadeMux I__927 (
            .O(N__4838),
            .I(N__4834));
    InMux I__926 (
            .O(N__4837),
            .I(N__4829));
    InMux I__925 (
            .O(N__4834),
            .I(N__4826));
    InMux I__924 (
            .O(N__4833),
            .I(N__4823));
    InMux I__923 (
            .O(N__4832),
            .I(N__4820));
    LocalMux I__922 (
            .O(N__4829),
            .I(N__4817));
    LocalMux I__921 (
            .O(N__4826),
            .I(\pc.program_counterZ0Z_1 ));
    LocalMux I__920 (
            .O(N__4823),
            .I(\pc.program_counterZ0Z_1 ));
    LocalMux I__919 (
            .O(N__4820),
            .I(\pc.program_counterZ0Z_1 ));
    Odrv12 I__918 (
            .O(N__4817),
            .I(\pc.program_counterZ0Z_1 ));
    ClkMux I__917 (
            .O(N__4808),
            .I(N__4700));
    ClkMux I__916 (
            .O(N__4807),
            .I(N__4700));
    ClkMux I__915 (
            .O(N__4806),
            .I(N__4700));
    ClkMux I__914 (
            .O(N__4805),
            .I(N__4700));
    ClkMux I__913 (
            .O(N__4804),
            .I(N__4700));
    ClkMux I__912 (
            .O(N__4803),
            .I(N__4700));
    ClkMux I__911 (
            .O(N__4802),
            .I(N__4700));
    ClkMux I__910 (
            .O(N__4801),
            .I(N__4700));
    ClkMux I__909 (
            .O(N__4800),
            .I(N__4700));
    ClkMux I__908 (
            .O(N__4799),
            .I(N__4700));
    ClkMux I__907 (
            .O(N__4798),
            .I(N__4700));
    ClkMux I__906 (
            .O(N__4797),
            .I(N__4700));
    ClkMux I__905 (
            .O(N__4796),
            .I(N__4700));
    ClkMux I__904 (
            .O(N__4795),
            .I(N__4700));
    ClkMux I__903 (
            .O(N__4794),
            .I(N__4700));
    ClkMux I__902 (
            .O(N__4793),
            .I(N__4700));
    ClkMux I__901 (
            .O(N__4792),
            .I(N__4700));
    ClkMux I__900 (
            .O(N__4791),
            .I(N__4700));
    ClkMux I__899 (
            .O(N__4790),
            .I(N__4700));
    ClkMux I__898 (
            .O(N__4789),
            .I(N__4700));
    ClkMux I__897 (
            .O(N__4788),
            .I(N__4700));
    ClkMux I__896 (
            .O(N__4787),
            .I(N__4700));
    ClkMux I__895 (
            .O(N__4786),
            .I(N__4700));
    ClkMux I__894 (
            .O(N__4785),
            .I(N__4700));
    ClkMux I__893 (
            .O(N__4784),
            .I(N__4700));
    ClkMux I__892 (
            .O(N__4783),
            .I(N__4700));
    ClkMux I__891 (
            .O(N__4782),
            .I(N__4700));
    ClkMux I__890 (
            .O(N__4781),
            .I(N__4700));
    ClkMux I__889 (
            .O(N__4780),
            .I(N__4700));
    ClkMux I__888 (
            .O(N__4779),
            .I(N__4700));
    ClkMux I__887 (
            .O(N__4778),
            .I(N__4700));
    ClkMux I__886 (
            .O(N__4777),
            .I(N__4700));
    ClkMux I__885 (
            .O(N__4776),
            .I(N__4700));
    ClkMux I__884 (
            .O(N__4775),
            .I(N__4700));
    ClkMux I__883 (
            .O(N__4774),
            .I(N__4700));
    ClkMux I__882 (
            .O(N__4773),
            .I(N__4700));
    GlobalMux I__881 (
            .O(N__4700),
            .I(N__4697));
    gio2CtrlBuf I__880 (
            .O(N__4697),
            .I(buf_clk_1_g));
    CascadeMux I__879 (
            .O(N__4694),
            .I(N__4687));
    InMux I__878 (
            .O(N__4693),
            .I(N__4681));
    InMux I__877 (
            .O(N__4692),
            .I(N__4681));
    InMux I__876 (
            .O(N__4691),
            .I(N__4678));
    InMux I__875 (
            .O(N__4690),
            .I(N__4673));
    InMux I__874 (
            .O(N__4687),
            .I(N__4673));
    CascadeMux I__873 (
            .O(N__4686),
            .I(N__4670));
    LocalMux I__872 (
            .O(N__4681),
            .I(N__4663));
    LocalMux I__871 (
            .O(N__4678),
            .I(N__4658));
    LocalMux I__870 (
            .O(N__4673),
            .I(N__4658));
    InMux I__869 (
            .O(N__4670),
            .I(N__4655));
    InMux I__868 (
            .O(N__4669),
            .I(N__4651));
    CascadeMux I__867 (
            .O(N__4668),
            .I(N__4648));
    InMux I__866 (
            .O(N__4667),
            .I(N__4645));
    CascadeMux I__865 (
            .O(N__4666),
            .I(N__4641));
    Span4Mux_h I__864 (
            .O(N__4663),
            .I(N__4632));
    Span4Mux_v I__863 (
            .O(N__4658),
            .I(N__4632));
    LocalMux I__862 (
            .O(N__4655),
            .I(N__4632));
    CascadeMux I__861 (
            .O(N__4654),
            .I(N__4629));
    LocalMux I__860 (
            .O(N__4651),
            .I(N__4626));
    InMux I__859 (
            .O(N__4648),
            .I(N__4623));
    LocalMux I__858 (
            .O(N__4645),
            .I(N__4620));
    InMux I__857 (
            .O(N__4644),
            .I(N__4615));
    InMux I__856 (
            .O(N__4641),
            .I(N__4615));
    InMux I__855 (
            .O(N__4640),
            .I(N__4610));
    InMux I__854 (
            .O(N__4639),
            .I(N__4610));
    Span4Mux_h I__853 (
            .O(N__4632),
            .I(N__4607));
    InMux I__852 (
            .O(N__4629),
            .I(N__4604));
    Odrv4 I__851 (
            .O(N__4626),
            .I(seq_T_2));
    LocalMux I__850 (
            .O(N__4623),
            .I(seq_T_2));
    Odrv12 I__849 (
            .O(N__4620),
            .I(seq_T_2));
    LocalMux I__848 (
            .O(N__4615),
            .I(seq_T_2));
    LocalMux I__847 (
            .O(N__4610),
            .I(seq_T_2));
    Odrv4 I__846 (
            .O(N__4607),
            .I(seq_T_2));
    LocalMux I__845 (
            .O(N__4604),
            .I(seq_T_2));
    InMux I__844 (
            .O(N__4589),
            .I(N__4584));
    InMux I__843 (
            .O(N__4588),
            .I(N__4581));
    InMux I__842 (
            .O(N__4587),
            .I(N__4574));
    LocalMux I__841 (
            .O(N__4584),
            .I(N__4571));
    LocalMux I__840 (
            .O(N__4581),
            .I(N__4568));
    InMux I__839 (
            .O(N__4580),
            .I(N__4563));
    InMux I__838 (
            .O(N__4579),
            .I(N__4563));
    InMux I__837 (
            .O(N__4578),
            .I(N__4558));
    InMux I__836 (
            .O(N__4577),
            .I(N__4558));
    LocalMux I__835 (
            .O(N__4574),
            .I(N__4555));
    Span4Mux_v I__834 (
            .O(N__4571),
            .I(N__4548));
    Span4Mux_v I__833 (
            .O(N__4568),
            .I(N__4548));
    LocalMux I__832 (
            .O(N__4563),
            .I(N__4548));
    LocalMux I__831 (
            .O(N__4558),
            .I(N__4544));
    Span4Mux_s2_v I__830 (
            .O(N__4555),
            .I(N__4536));
    Span4Mux_h I__829 (
            .O(N__4548),
            .I(N__4533));
    InMux I__828 (
            .O(N__4547),
            .I(N__4530));
    Span4Mux_h I__827 (
            .O(N__4544),
            .I(N__4527));
    InMux I__826 (
            .O(N__4543),
            .I(N__4522));
    InMux I__825 (
            .O(N__4542),
            .I(N__4522));
    InMux I__824 (
            .O(N__4541),
            .I(N__4515));
    InMux I__823 (
            .O(N__4540),
            .I(N__4515));
    InMux I__822 (
            .O(N__4539),
            .I(N__4515));
    Odrv4 I__821 (
            .O(N__4536),
            .I(seq_PC_LD_0_0));
    Odrv4 I__820 (
            .O(N__4533),
            .I(seq_PC_LD_0_0));
    LocalMux I__819 (
            .O(N__4530),
            .I(seq_PC_LD_0_0));
    Odrv4 I__818 (
            .O(N__4527),
            .I(seq_PC_LD_0_0));
    LocalMux I__817 (
            .O(N__4522),
            .I(seq_PC_LD_0_0));
    LocalMux I__816 (
            .O(N__4515),
            .I(seq_PC_LD_0_0));
    InMux I__815 (
            .O(N__4502),
            .I(N__4498));
    InMux I__814 (
            .O(N__4501),
            .I(N__4494));
    LocalMux I__813 (
            .O(N__4498),
            .I(N__4489));
    InMux I__812 (
            .O(N__4497),
            .I(N__4486));
    LocalMux I__811 (
            .O(N__4494),
            .I(N__4482));
    InMux I__810 (
            .O(N__4493),
            .I(N__4479));
    InMux I__809 (
            .O(N__4492),
            .I(N__4476));
    Span4Mux_v I__808 (
            .O(N__4489),
            .I(N__4473));
    LocalMux I__807 (
            .O(N__4486),
            .I(N__4470));
    InMux I__806 (
            .O(N__4485),
            .I(N__4467));
    Span4Mux_v I__805 (
            .O(N__4482),
            .I(N__4462));
    LocalMux I__804 (
            .O(N__4479),
            .I(N__4462));
    LocalMux I__803 (
            .O(N__4476),
            .I(N__4459));
    Span4Mux_v I__802 (
            .O(N__4473),
            .I(N__4454));
    Span4Mux_v I__801 (
            .O(N__4470),
            .I(N__4447));
    LocalMux I__800 (
            .O(N__4467),
            .I(N__4447));
    Span4Mux_h I__799 (
            .O(N__4462),
            .I(N__4447));
    Span4Mux_h I__798 (
            .O(N__4459),
            .I(N__4444));
    InMux I__797 (
            .O(N__4458),
            .I(N__4439));
    InMux I__796 (
            .O(N__4457),
            .I(N__4439));
    Odrv4 I__795 (
            .O(N__4454),
            .I(seq_MAR_LD_2));
    Odrv4 I__794 (
            .O(N__4447),
            .I(seq_MAR_LD_2));
    Odrv4 I__793 (
            .O(N__4444),
            .I(seq_MAR_LD_2));
    LocalMux I__792 (
            .O(N__4439),
            .I(seq_MAR_LD_2));
    CascadeMux I__791 (
            .O(N__4430),
            .I(N__4427));
    InMux I__790 (
            .O(N__4427),
            .I(N__4424));
    LocalMux I__789 (
            .O(N__4424),
            .I(N__4421));
    Odrv4 I__788 (
            .O(N__4421),
            .I(\seq.gZ0Z2 ));
    InMux I__787 (
            .O(N__4418),
            .I(N__4414));
    InMux I__786 (
            .O(N__4417),
            .I(N__4408));
    LocalMux I__785 (
            .O(N__4414),
            .I(N__4405));
    InMux I__784 (
            .O(N__4413),
            .I(N__4402));
    InMux I__783 (
            .O(N__4412),
            .I(N__4397));
    InMux I__782 (
            .O(N__4411),
            .I(N__4397));
    LocalMux I__781 (
            .O(N__4408),
            .I(ir_out_5));
    Odrv4 I__780 (
            .O(N__4405),
            .I(ir_out_5));
    LocalMux I__779 (
            .O(N__4402),
            .I(ir_out_5));
    LocalMux I__778 (
            .O(N__4397),
            .I(ir_out_5));
    InMux I__777 (
            .O(N__4388),
            .I(N__4384));
    InMux I__776 (
            .O(N__4387),
            .I(N__4380));
    LocalMux I__775 (
            .O(N__4384),
            .I(N__4377));
    InMux I__774 (
            .O(N__4383),
            .I(N__4374));
    LocalMux I__773 (
            .O(N__4380),
            .I(N__4369));
    Span4Mux_h I__772 (
            .O(N__4377),
            .I(N__4369));
    LocalMux I__771 (
            .O(N__4374),
            .I(N__4366));
    Span4Mux_v I__770 (
            .O(N__4369),
            .I(N__4363));
    Odrv4 I__769 (
            .O(N__4366),
            .I(bus_7));
    Odrv4 I__768 (
            .O(N__4363),
            .I(bus_7));
    InMux I__767 (
            .O(N__4358),
            .I(N__4355));
    LocalMux I__766 (
            .O(N__4355),
            .I(N__4352));
    Span4Mux_s2_v I__765 (
            .O(N__4352),
            .I(N__4348));
    InMux I__764 (
            .O(N__4351),
            .I(N__4345));
    Odrv4 I__763 (
            .O(N__4348),
            .I(N_5_0));
    LocalMux I__762 (
            .O(N__4345),
            .I(N_5_0));
    CascadeMux I__761 (
            .O(N__4340),
            .I(N_1_0_cascade_));
    InMux I__760 (
            .O(N__4337),
            .I(N__4334));
    LocalMux I__759 (
            .O(N__4334),
            .I(N__4331));
    Span4Mux_v I__758 (
            .O(N__4331),
            .I(N__4328));
    Span4Mux_v I__757 (
            .O(N__4328),
            .I(N__4325));
    Odrv4 I__756 (
            .O(N__4325),
            .I(seq_un1_HLT_0));
    InMux I__755 (
            .O(N__4322),
            .I(N__4319));
    LocalMux I__754 (
            .O(N__4319),
            .I(\seq.un1_HLT_1_reti ));
    InMux I__753 (
            .O(N__4316),
            .I(N__4313));
    LocalMux I__752 (
            .O(N__4313),
            .I(N__4310));
    Span4Mux_s3_h I__751 (
            .O(N__4310),
            .I(N__4305));
    InMux I__750 (
            .O(N__4309),
            .I(N__4302));
    InMux I__749 (
            .O(N__4308),
            .I(N__4299));
    Odrv4 I__748 (
            .O(N__4305),
            .I(N_2_0));
    LocalMux I__747 (
            .O(N__4302),
            .I(N_2_0));
    LocalMux I__746 (
            .O(N__4299),
            .I(N_2_0));
    CascadeMux I__745 (
            .O(N__4292),
            .I(N__4289));
    InMux I__744 (
            .O(N__4289),
            .I(N__4286));
    LocalMux I__743 (
            .O(N__4286),
            .I(N__4283));
    Span4Mux_v I__742 (
            .O(N__4283),
            .I(N__4280));
    Odrv4 I__741 (
            .O(N__4280),
            .I(\seq.un1_HLT_1 ));
    CascadeMux I__740 (
            .O(N__4277),
            .I(bus_1_cascade_));
    InMux I__739 (
            .O(N__4274),
            .I(N__4268));
    InMux I__738 (
            .O(N__4273),
            .I(N__4264));
    InMux I__737 (
            .O(N__4272),
            .I(N__4259));
    InMux I__736 (
            .O(N__4271),
            .I(N__4259));
    LocalMux I__735 (
            .O(N__4268),
            .I(N__4256));
    InMux I__734 (
            .O(N__4267),
            .I(N__4253));
    LocalMux I__733 (
            .O(N__4264),
            .I(N__4243));
    LocalMux I__732 (
            .O(N__4259),
            .I(N__4243));
    Span4Mux_v I__731 (
            .O(N__4256),
            .I(N__4238));
    LocalMux I__730 (
            .O(N__4253),
            .I(N__4238));
    InMux I__729 (
            .O(N__4252),
            .I(N__4233));
    InMux I__728 (
            .O(N__4251),
            .I(N__4233));
    InMux I__727 (
            .O(N__4250),
            .I(N__4228));
    InMux I__726 (
            .O(N__4249),
            .I(N__4228));
    InMux I__725 (
            .O(N__4248),
            .I(N__4225));
    Odrv4 I__724 (
            .O(N__4243),
            .I(seq_D_6));
    Odrv4 I__723 (
            .O(N__4238),
            .I(seq_D_6));
    LocalMux I__722 (
            .O(N__4233),
            .I(seq_D_6));
    LocalMux I__721 (
            .O(N__4228),
            .I(seq_D_6));
    LocalMux I__720 (
            .O(N__4225),
            .I(seq_D_6));
    InMux I__719 (
            .O(N__4214),
            .I(N__4210));
    InMux I__718 (
            .O(N__4213),
            .I(N__4207));
    LocalMux I__717 (
            .O(N__4210),
            .I(N__4198));
    LocalMux I__716 (
            .O(N__4207),
            .I(N__4198));
    InMux I__715 (
            .O(N__4206),
            .I(N__4195));
    InMux I__714 (
            .O(N__4205),
            .I(N__4191));
    InMux I__713 (
            .O(N__4204),
            .I(N__4188));
    InMux I__712 (
            .O(N__4203),
            .I(N__4185));
    Span4Mux_h I__711 (
            .O(N__4198),
            .I(N__4180));
    LocalMux I__710 (
            .O(N__4195),
            .I(N__4176));
    InMux I__709 (
            .O(N__4194),
            .I(N__4173));
    LocalMux I__708 (
            .O(N__4191),
            .I(N__4166));
    LocalMux I__707 (
            .O(N__4188),
            .I(N__4166));
    LocalMux I__706 (
            .O(N__4185),
            .I(N__4166));
    InMux I__705 (
            .O(N__4184),
            .I(N__4161));
    InMux I__704 (
            .O(N__4183),
            .I(N__4161));
    Span4Mux_v I__703 (
            .O(N__4180),
            .I(N__4158));
    InMux I__702 (
            .O(N__4179),
            .I(N__4155));
    Span4Mux_h I__701 (
            .O(N__4176),
            .I(N__4150));
    LocalMux I__700 (
            .O(N__4173),
            .I(N__4150));
    Span4Mux_v I__699 (
            .O(N__4166),
            .I(N__4147));
    LocalMux I__698 (
            .O(N__4161),
            .I(T_0_fast_RNILB791_2));
    Odrv4 I__697 (
            .O(N__4158),
            .I(T_0_fast_RNILB791_2));
    LocalMux I__696 (
            .O(N__4155),
            .I(T_0_fast_RNILB791_2));
    Odrv4 I__695 (
            .O(N__4150),
            .I(T_0_fast_RNILB791_2));
    Odrv4 I__694 (
            .O(N__4147),
            .I(T_0_fast_RNILB791_2));
    CascadeMux I__693 (
            .O(N__4136),
            .I(N__4132));
    InMux I__692 (
            .O(N__4135),
            .I(N__4129));
    InMux I__691 (
            .O(N__4132),
            .I(N__4126));
    LocalMux I__690 (
            .O(N__4129),
            .I(AR_out_1));
    LocalMux I__689 (
            .O(N__4126),
            .I(AR_out_1));
    CascadeMux I__688 (
            .O(N__4121),
            .I(ALU_main_N_44_0_cascade_));
    InMux I__687 (
            .O(N__4118),
            .I(N__4112));
    InMux I__686 (
            .O(N__4117),
            .I(N__4112));
    LocalMux I__685 (
            .O(N__4112),
            .I(un1_A_cry_2_c_RNI1TTO2));
    InMux I__684 (
            .O(N__4109),
            .I(N__4106));
    LocalMux I__683 (
            .O(N__4106),
            .I(N__4103));
    Odrv4 I__682 (
            .O(N__4103),
            .I(\pc.N_10_i ));
    InMux I__681 (
            .O(N__4100),
            .I(N__4097));
    LocalMux I__680 (
            .O(N__4097),
            .I(N__4094));
    Span12Mux_s4_v I__679 (
            .O(N__4094),
            .I(N__4091));
    Odrv12 I__678 (
            .O(N__4091),
            .I(\pc.G_10_0_1_1 ));
    InMux I__677 (
            .O(N__4088),
            .I(N__4085));
    LocalMux I__676 (
            .O(N__4085),
            .I(N__4082));
    Odrv4 I__675 (
            .O(N__4082),
            .I(\pc.G_10_0_1 ));
    CascadeMux I__674 (
            .O(N__4079),
            .I(N__4076));
    InMux I__673 (
            .O(N__4076),
            .I(N__4073));
    LocalMux I__672 (
            .O(N__4073),
            .I(ALU_main_N_44_1));
    InMux I__671 (
            .O(N__4070),
            .I(N__4067));
    LocalMux I__670 (
            .O(N__4067),
            .I(N__4064));
    Odrv12 I__669 (
            .O(N__4064),
            .I(\pc.un1_inc_0_0 ));
    InMux I__668 (
            .O(N__4061),
            .I(N__4058));
    LocalMux I__667 (
            .O(N__4058),
            .I(N__4055));
    Span4Mux_v I__666 (
            .O(N__4055),
            .I(N__4052));
    Odrv4 I__665 (
            .O(N__4052),
            .I(\pc.out_1_iv_1_1 ));
    CascadeMux I__664 (
            .O(N__4049),
            .I(N__4046));
    InMux I__663 (
            .O(N__4046),
            .I(N__4043));
    LocalMux I__662 (
            .O(N__4043),
            .I(N__4040));
    Span4Mux_v I__661 (
            .O(N__4040),
            .I(N__4037));
    Span4Mux_h I__660 (
            .O(N__4037),
            .I(N__4034));
    Odrv4 I__659 (
            .O(N__4034),
            .I(mem_data_2_7_0__N_16_0));
    InMux I__658 (
            .O(N__4031),
            .I(N__4028));
    LocalMux I__657 (
            .O(N__4028),
            .I(N__4025));
    Span4Mux_h I__656 (
            .O(N__4025),
            .I(N__4022));
    Odrv4 I__655 (
            .O(N__4022),
            .I(\pc.g0_rn_1 ));
    CascadeMux I__654 (
            .O(N__4019),
            .I(\pc.g0_sn_cascade_ ));
    InMux I__653 (
            .O(N__4016),
            .I(N__4013));
    LocalMux I__652 (
            .O(N__4013),
            .I(alu_out_m_0_3));
    InMux I__651 (
            .O(N__4010),
            .I(N__4006));
    InMux I__650 (
            .O(N__4009),
            .I(N__4003));
    LocalMux I__649 (
            .O(N__4006),
            .I(N__4000));
    LocalMux I__648 (
            .O(N__4003),
            .I(N__3997));
    Span4Mux_v I__647 (
            .O(N__4000),
            .I(N__3992));
    Span4Mux_s3_h I__646 (
            .O(N__3997),
            .I(N__3992));
    Odrv4 I__645 (
            .O(N__3992),
            .I(\pc.program_counterZ0Z_3 ));
    InMux I__644 (
            .O(N__3989),
            .I(N__3986));
    LocalMux I__643 (
            .O(N__3986),
            .I(N__3982));
    InMux I__642 (
            .O(N__3985),
            .I(N__3979));
    Span4Mux_h I__641 (
            .O(N__3982),
            .I(N__3976));
    LocalMux I__640 (
            .O(N__3979),
            .I(seq_un1_AR_OE_0_0));
    Odrv4 I__639 (
            .O(N__3976),
            .I(seq_un1_AR_OE_0_0));
    InMux I__638 (
            .O(N__3971),
            .I(N__3968));
    LocalMux I__637 (
            .O(N__3968),
            .I(N__3960));
    InMux I__636 (
            .O(N__3967),
            .I(N__3955));
    InMux I__635 (
            .O(N__3966),
            .I(N__3955));
    CascadeMux I__634 (
            .O(N__3965),
            .I(N__3952));
    InMux I__633 (
            .O(N__3964),
            .I(N__3949));
    InMux I__632 (
            .O(N__3963),
            .I(N__3946));
    Span4Mux_v I__631 (
            .O(N__3960),
            .I(N__3943));
    LocalMux I__630 (
            .O(N__3955),
            .I(N__3940));
    InMux I__629 (
            .O(N__3952),
            .I(N__3937));
    LocalMux I__628 (
            .O(N__3949),
            .I(ir_out_6));
    LocalMux I__627 (
            .O(N__3946),
            .I(ir_out_6));
    Odrv4 I__626 (
            .O(N__3943),
            .I(ir_out_6));
    Odrv12 I__625 (
            .O(N__3940),
            .I(ir_out_6));
    LocalMux I__624 (
            .O(N__3937),
            .I(ir_out_6));
    InMux I__623 (
            .O(N__3926),
            .I(N__3922));
    CascadeMux I__622 (
            .O(N__3925),
            .I(N__3919));
    LocalMux I__621 (
            .O(N__3922),
            .I(N__3916));
    InMux I__620 (
            .O(N__3919),
            .I(N__3913));
    Span4Mux_s1_v I__619 (
            .O(N__3916),
            .I(N__3909));
    LocalMux I__618 (
            .O(N__3913),
            .I(N__3906));
    InMux I__617 (
            .O(N__3912),
            .I(N__3903));
    Span4Mux_v I__616 (
            .O(N__3909),
            .I(N__3900));
    Span4Mux_h I__615 (
            .O(N__3906),
            .I(N__3897));
    LocalMux I__614 (
            .O(N__3903),
            .I(\AR.ff4.AR_out_3 ));
    Odrv4 I__613 (
            .O(N__3900),
            .I(\AR.ff4.AR_out_3 ));
    Odrv4 I__612 (
            .O(N__3897),
            .I(\AR.ff4.AR_out_3 ));
    InMux I__611 (
            .O(N__3890),
            .I(N__3885));
    InMux I__610 (
            .O(N__3889),
            .I(N__3882));
    InMux I__609 (
            .O(N__3888),
            .I(N__3879));
    LocalMux I__608 (
            .O(N__3885),
            .I(N__3876));
    LocalMux I__607 (
            .O(N__3882),
            .I(N__3872));
    LocalMux I__606 (
            .O(N__3879),
            .I(N__3869));
    Span4Mux_v I__605 (
            .O(N__3876),
            .I(N__3866));
    InMux I__604 (
            .O(N__3875),
            .I(N__3863));
    Span4Mux_h I__603 (
            .O(N__3872),
            .I(N__3860));
    Span4Mux_s2_h I__602 (
            .O(N__3869),
            .I(N__3857));
    Odrv4 I__601 (
            .O(N__3866),
            .I(ir_out_3));
    LocalMux I__600 (
            .O(N__3863),
            .I(ir_out_3));
    Odrv4 I__599 (
            .O(N__3860),
            .I(ir_out_3));
    Odrv4 I__598 (
            .O(N__3857),
            .I(ir_out_3));
    InMux I__597 (
            .O(N__3848),
            .I(N__3845));
    LocalMux I__596 (
            .O(N__3845),
            .I(\pc.tbuf.g0_0_1_0 ));
    CascadeMux I__595 (
            .O(N__3842),
            .I(AR_out_m_3_cascade_));
    InMux I__594 (
            .O(N__3839),
            .I(N__3836));
    LocalMux I__593 (
            .O(N__3836),
            .I(\pc.g0_0 ));
    CascadeMux I__592 (
            .O(N__3833),
            .I(N__3830));
    InMux I__591 (
            .O(N__3830),
            .I(N__3827));
    LocalMux I__590 (
            .O(N__3827),
            .I(\ALU_main.un1_A_axb_2_l_ofxZ0 ));
    InMux I__589 (
            .O(N__3824),
            .I(N__3821));
    LocalMux I__588 (
            .O(N__3821),
            .I(N__3817));
    InMux I__587 (
            .O(N__3820),
            .I(N__3814));
    Odrv4 I__586 (
            .O(N__3817),
            .I(un1_A_cry_1_c_RNITKPO2));
    LocalMux I__585 (
            .O(N__3814),
            .I(un1_A_cry_1_c_RNITKPO2));
    InMux I__584 (
            .O(N__3809),
            .I(\ALU_main.un1_A_cry_1 ));
    InMux I__583 (
            .O(N__3806),
            .I(\ALU_main.un1_A_cry_2 ));
    InMux I__582 (
            .O(N__3803),
            .I(\ALU_main.un1_A_cry_3 ));
    InMux I__581 (
            .O(N__3800),
            .I(\ALU_main.un1_A_cry_4 ));
    InMux I__580 (
            .O(N__3797),
            .I(\ALU_main.un1_A_cry_5 ));
    InMux I__579 (
            .O(N__3794),
            .I(bfn_4_13_0_));
    InMux I__578 (
            .O(N__3791),
            .I(N__3788));
    LocalMux I__577 (
            .O(N__3788),
            .I(N__3785));
    Span4Mux_s3_h I__576 (
            .O(N__3785),
            .I(N__3782));
    Odrv4 I__575 (
            .O(N__3782),
            .I(\ALU_main.un1_A_cry_6_c_RNIP89EZ0Z2 ));
    InMux I__574 (
            .O(N__3779),
            .I(N__3776));
    LocalMux I__573 (
            .O(N__3776),
            .I(\ALU_main.un1_A_cry_5_c_RNIDLAPZ0Z2 ));
    InMux I__572 (
            .O(N__3773),
            .I(N__3770));
    LocalMux I__571 (
            .O(N__3770),
            .I(N__3766));
    InMux I__570 (
            .O(N__3769),
            .I(N__3763));
    Span4Mux_h I__569 (
            .O(N__3766),
            .I(N__3760));
    LocalMux I__568 (
            .O(N__3763),
            .I(N__3757));
    Odrv4 I__567 (
            .O(N__3760),
            .I(N_30));
    Odrv4 I__566 (
            .O(N__3757),
            .I(N_30));
    CascadeMux I__565 (
            .O(N__3752),
            .I(\pc.G_10_0_1_0_cascade_ ));
    InMux I__564 (
            .O(N__3749),
            .I(N__3746));
    LocalMux I__563 (
            .O(N__3746),
            .I(N__3743));
    Odrv4 I__562 (
            .O(N__3743),
            .I(\pc.G_10_0_sx ));
    CascadeMux I__561 (
            .O(N__3740),
            .I(N__3737));
    InMux I__560 (
            .O(N__3737),
            .I(N__3734));
    LocalMux I__559 (
            .O(N__3734),
            .I(\pc.G_10_0_5_1 ));
    InMux I__558 (
            .O(N__3731),
            .I(N__3728));
    LocalMux I__557 (
            .O(N__3728),
            .I(N__3725));
    Odrv4 I__556 (
            .O(N__3725),
            .I(ALU_main_N_43_0));
    CascadeMux I__555 (
            .O(N__3722),
            .I(N__3719));
    InMux I__554 (
            .O(N__3719),
            .I(N__3715));
    InMux I__553 (
            .O(N__3718),
            .I(N__3712));
    LocalMux I__552 (
            .O(N__3715),
            .I(N__3708));
    LocalMux I__551 (
            .O(N__3712),
            .I(N__3705));
    InMux I__550 (
            .O(N__3711),
            .I(N__3701));
    Span4Mux_v I__549 (
            .O(N__3708),
            .I(N__3695));
    Span4Mux_v I__548 (
            .O(N__3705),
            .I(N__3695));
    InMux I__547 (
            .O(N__3704),
            .I(N__3692));
    LocalMux I__546 (
            .O(N__3701),
            .I(N__3689));
    InMux I__545 (
            .O(N__3700),
            .I(N__3686));
    Span4Mux_h I__544 (
            .O(N__3695),
            .I(N__3681));
    LocalMux I__543 (
            .O(N__3692),
            .I(N__3681));
    Span4Mux_s3_h I__542 (
            .O(N__3689),
            .I(N__3678));
    LocalMux I__541 (
            .O(N__3686),
            .I(\pc.program_counterZ0Z_2 ));
    Odrv4 I__540 (
            .O(N__3681),
            .I(\pc.program_counterZ0Z_2 ));
    Odrv4 I__539 (
            .O(N__3678),
            .I(\pc.program_counterZ0Z_2 ));
    InMux I__538 (
            .O(N__3671),
            .I(N__3667));
    InMux I__537 (
            .O(N__3670),
            .I(N__3663));
    LocalMux I__536 (
            .O(N__3667),
            .I(N__3659));
    InMux I__535 (
            .O(N__3666),
            .I(N__3656));
    LocalMux I__534 (
            .O(N__3663),
            .I(N__3653));
    InMux I__533 (
            .O(N__3662),
            .I(N__3650));
    Span4Mux_h I__532 (
            .O(N__3659),
            .I(N__3645));
    LocalMux I__531 (
            .O(N__3656),
            .I(N__3645));
    Span4Mux_v I__530 (
            .O(N__3653),
            .I(N__3636));
    LocalMux I__529 (
            .O(N__3650),
            .I(N__3636));
    Span4Mux_v I__528 (
            .O(N__3645),
            .I(N__3636));
    InMux I__527 (
            .O(N__3644),
            .I(N__3631));
    InMux I__526 (
            .O(N__3643),
            .I(N__3631));
    Odrv4 I__525 (
            .O(N__3636),
            .I(\pc.program_counterZ0Z_0 ));
    LocalMux I__524 (
            .O(N__3631),
            .I(\pc.program_counterZ0Z_0 ));
    CascadeMux I__523 (
            .O(N__3626),
            .I(N__3623));
    InMux I__522 (
            .O(N__3623),
            .I(N__3619));
    InMux I__521 (
            .O(N__3622),
            .I(N__3616));
    LocalMux I__520 (
            .O(N__3619),
            .I(N__3611));
    LocalMux I__519 (
            .O(N__3616),
            .I(N__3611));
    Odrv4 I__518 (
            .O(N__3611),
            .I(seq_S0_0_i));
    InMux I__517 (
            .O(N__3608),
            .I(\ALU_main.un1_A_cry_0_c_THRU_CO ));
    InMux I__516 (
            .O(N__3605),
            .I(\ALU_main.un1_A_cry_0 ));
    CascadeMux I__515 (
            .O(N__3602),
            .I(IR_OE_1_cascade_));
    InMux I__514 (
            .O(N__3599),
            .I(N__3593));
    InMux I__513 (
            .O(N__3598),
            .I(N__3593));
    LocalMux I__512 (
            .O(N__3593),
            .I(\pc.un1_inc_0 ));
    CascadeMux I__511 (
            .O(N__3590),
            .I(N__3587));
    InMux I__510 (
            .O(N__3587),
            .I(N__3584));
    LocalMux I__509 (
            .O(N__3584),
            .I(N__3581));
    Odrv12 I__508 (
            .O(N__3581),
            .I(\pc.G_12_i_a3_2_3 ));
    InMux I__507 (
            .O(N__3578),
            .I(N__3575));
    LocalMux I__506 (
            .O(N__3575),
            .I(\pc.G_12_i_a3_2_1 ));
    CascadeMux I__505 (
            .O(N__3572),
            .I(\seq.counter.T8_1_cascade_ ));
    CascadeMux I__504 (
            .O(N__3569),
            .I(N__3566));
    InMux I__503 (
            .O(N__3566),
            .I(N__3563));
    LocalMux I__502 (
            .O(N__3563),
            .I(\pc.g1_0 ));
    InMux I__501 (
            .O(N__3560),
            .I(N__3557));
    LocalMux I__500 (
            .O(N__3557),
            .I(N__3554));
    Span4Mux_s3_h I__499 (
            .O(N__3554),
            .I(N__3551));
    Odrv4 I__498 (
            .O(N__3551),
            .I(\pc.N_188_0 ));
    CascadeMux I__497 (
            .O(N__3548),
            .I(N__3542));
    CascadeMux I__496 (
            .O(N__3547),
            .I(N__3538));
    InMux I__495 (
            .O(N__3546),
            .I(N__3534));
    InMux I__494 (
            .O(N__3545),
            .I(N__3527));
    InMux I__493 (
            .O(N__3542),
            .I(N__3527));
    InMux I__492 (
            .O(N__3541),
            .I(N__3527));
    InMux I__491 (
            .O(N__3538),
            .I(N__3524));
    CascadeMux I__490 (
            .O(N__3537),
            .I(N__3520));
    LocalMux I__489 (
            .O(N__3534),
            .I(N__3517));
    LocalMux I__488 (
            .O(N__3527),
            .I(N__3511));
    LocalMux I__487 (
            .O(N__3524),
            .I(N__3508));
    InMux I__486 (
            .O(N__3523),
            .I(N__3503));
    InMux I__485 (
            .O(N__3520),
            .I(N__3503));
    Span4Mux_v I__484 (
            .O(N__3517),
            .I(N__3500));
    InMux I__483 (
            .O(N__3516),
            .I(N__3493));
    InMux I__482 (
            .O(N__3515),
            .I(N__3493));
    InMux I__481 (
            .O(N__3514),
            .I(N__3493));
    Span4Mux_v I__480 (
            .O(N__3511),
            .I(N__3486));
    Span4Mux_v I__479 (
            .O(N__3508),
            .I(N__3486));
    LocalMux I__478 (
            .O(N__3503),
            .I(N__3486));
    Odrv4 I__477 (
            .O(N__3500),
            .I(seq_T_0));
    LocalMux I__476 (
            .O(N__3493),
            .I(seq_T_0));
    Odrv4 I__475 (
            .O(N__3486),
            .I(seq_T_0));
    CascadeMux I__474 (
            .O(N__3479),
            .I(g0_0_1_cascade_));
    InMux I__473 (
            .O(N__3476),
            .I(N__3473));
    LocalMux I__472 (
            .O(N__3473),
            .I(N__3470));
    Odrv12 I__471 (
            .O(N__3470),
            .I(\seq.counter.un7_ACC_LD_0 ));
    InMux I__470 (
            .O(N__3467),
            .I(N__3464));
    LocalMux I__469 (
            .O(N__3464),
            .I(\seq.un1_ALU_en_0Z0Z_1 ));
    CascadeMux I__468 (
            .O(N__3461),
            .I(\seq.counter.un7_ACC_LD_0_cascade_ ));
    CascadeMux I__467 (
            .O(N__3458),
            .I(IR_OE_2_cascade_));
    InMux I__466 (
            .O(N__3455),
            .I(N__3452));
    LocalMux I__465 (
            .O(N__3452),
            .I(N__3449));
    Odrv4 I__464 (
            .O(N__3449),
            .I(bus_2));
    InMux I__463 (
            .O(N__3446),
            .I(N__3443));
    LocalMux I__462 (
            .O(N__3443),
            .I(N__3440));
    Span4Mux_h I__461 (
            .O(N__3440),
            .I(N__3437));
    Odrv4 I__460 (
            .O(N__3437),
            .I(\seq.g2Z0Z_0 ));
    InMux I__459 (
            .O(N__3434),
            .I(N__3429));
    CascadeMux I__458 (
            .O(N__3433),
            .I(N__3425));
    CascadeMux I__457 (
            .O(N__3432),
            .I(N__3421));
    LocalMux I__456 (
            .O(N__3429),
            .I(N__3418));
    InMux I__455 (
            .O(N__3428),
            .I(N__3413));
    InMux I__454 (
            .O(N__3425),
            .I(N__3413));
    CascadeMux I__453 (
            .O(N__3424),
            .I(N__3410));
    InMux I__452 (
            .O(N__3421),
            .I(N__3406));
    Span4Mux_s1_h I__451 (
            .O(N__3418),
            .I(N__3401));
    LocalMux I__450 (
            .O(N__3413),
            .I(N__3401));
    InMux I__449 (
            .O(N__3410),
            .I(N__3398));
    InMux I__448 (
            .O(N__3409),
            .I(N__3395));
    LocalMux I__447 (
            .O(N__3406),
            .I(ir_out_fast_7));
    Odrv4 I__446 (
            .O(N__3401),
            .I(ir_out_fast_7));
    LocalMux I__445 (
            .O(N__3398),
            .I(ir_out_fast_7));
    LocalMux I__444 (
            .O(N__3395),
            .I(ir_out_fast_7));
    InMux I__443 (
            .O(N__3386),
            .I(N__3383));
    LocalMux I__442 (
            .O(N__3383),
            .I(N__3380));
    Odrv4 I__441 (
            .O(N__3380),
            .I(\seq.S0_0_i_N_3LZ0Z3 ));
    InMux I__440 (
            .O(N__3377),
            .I(N__3371));
    InMux I__439 (
            .O(N__3376),
            .I(N__3366));
    InMux I__438 (
            .O(N__3375),
            .I(N__3366));
    InMux I__437 (
            .O(N__3374),
            .I(N__3363));
    LocalMux I__436 (
            .O(N__3371),
            .I(ir_out_i_2_6));
    LocalMux I__435 (
            .O(N__3366),
            .I(ir_out_i_2_6));
    LocalMux I__434 (
            .O(N__3363),
            .I(ir_out_i_2_6));
    InMux I__433 (
            .O(N__3356),
            .I(N__3352));
    CascadeMux I__432 (
            .O(N__3355),
            .I(N__3348));
    LocalMux I__431 (
            .O(N__3352),
            .I(N__3345));
    InMux I__430 (
            .O(N__3351),
            .I(N__3340));
    InMux I__429 (
            .O(N__3348),
            .I(N__3340));
    Odrv4 I__428 (
            .O(N__3345),
            .I(\seq.counter.T_fast_2 ));
    LocalMux I__427 (
            .O(N__3340),
            .I(\seq.counter.T_fast_2 ));
    InMux I__426 (
            .O(N__3335),
            .I(N__3332));
    LocalMux I__425 (
            .O(N__3332),
            .I(N__3329));
    Span4Mux_v I__424 (
            .O(N__3329),
            .I(N__3324));
    InMux I__423 (
            .O(N__3328),
            .I(N__3319));
    InMux I__422 (
            .O(N__3327),
            .I(N__3319));
    Odrv4 I__421 (
            .O(N__3324),
            .I(seq_un1_IR_OE_4_1));
    LocalMux I__420 (
            .O(N__3319),
            .I(seq_un1_IR_OE_4_1));
    CascadeMux I__419 (
            .O(N__3314),
            .I(\seq.B_LD_0_2_tz_cascade_ ));
    InMux I__418 (
            .O(N__3311),
            .I(N__3308));
    LocalMux I__417 (
            .O(N__3308),
            .I(N__3305));
    Odrv4 I__416 (
            .O(N__3305),
            .I(\seq.counter.T_RNIR83I4_0Z0Z_3 ));
    InMux I__415 (
            .O(N__3302),
            .I(N__3298));
    InMux I__414 (
            .O(N__3301),
            .I(N__3292));
    LocalMux I__413 (
            .O(N__3298),
            .I(N__3289));
    InMux I__412 (
            .O(N__3297),
            .I(N__3286));
    InMux I__411 (
            .O(N__3296),
            .I(N__3281));
    InMux I__410 (
            .O(N__3295),
            .I(N__3281));
    LocalMux I__409 (
            .O(N__3292),
            .I(IR_ff6_q_0_fast));
    Odrv12 I__408 (
            .O(N__3289),
            .I(IR_ff6_q_0_fast));
    LocalMux I__407 (
            .O(N__3286),
            .I(IR_ff6_q_0_fast));
    LocalMux I__406 (
            .O(N__3281),
            .I(IR_ff6_q_0_fast));
    InMux I__405 (
            .O(N__3272),
            .I(N__3269));
    LocalMux I__404 (
            .O(N__3269),
            .I(N__3262));
    InMux I__403 (
            .O(N__3268),
            .I(N__3255));
    InMux I__402 (
            .O(N__3267),
            .I(N__3255));
    InMux I__401 (
            .O(N__3266),
            .I(N__3255));
    InMux I__400 (
            .O(N__3265),
            .I(N__3252));
    Odrv4 I__399 (
            .O(N__3262),
            .I(IR_ff7_q_ret_1_fast));
    LocalMux I__398 (
            .O(N__3255),
            .I(IR_ff7_q_ret_1_fast));
    LocalMux I__397 (
            .O(N__3252),
            .I(IR_ff7_q_ret_1_fast));
    CascadeMux I__396 (
            .O(N__3245),
            .I(\seq.counter.T_0_fast_RNIP4D21Z0Z_2_cascade_ ));
    CascadeMux I__395 (
            .O(N__3242),
            .I(T_0_fast_RNILB791_2_cascade_));
    InMux I__394 (
            .O(N__3239),
            .I(N__3236));
    LocalMux I__393 (
            .O(N__3236),
            .I(N__3233));
    Span4Mux_s2_h I__392 (
            .O(N__3233),
            .I(N__3230));
    Odrv4 I__391 (
            .O(N__3230),
            .I(\pc.G_12_i_0 ));
    CascadeMux I__390 (
            .O(N__3227),
            .I(\seq.counter.T_0_fast_RNIG89VZ0Z_2_cascade_ ));
    InMux I__389 (
            .O(N__3224),
            .I(N__3221));
    LocalMux I__388 (
            .O(N__3221),
            .I(N__3218));
    Odrv4 I__387 (
            .O(N__3218),
            .I(bus_6));
    CascadeMux I__386 (
            .O(N__3215),
            .I(N__3212));
    InMux I__385 (
            .O(N__3212),
            .I(N__3207));
    InMux I__384 (
            .O(N__3211),
            .I(N__3202));
    InMux I__383 (
            .O(N__3210),
            .I(N__3202));
    LocalMux I__382 (
            .O(N__3207),
            .I(ir_out_fast_4));
    LocalMux I__381 (
            .O(N__3202),
            .I(ir_out_fast_4));
    CascadeMux I__380 (
            .O(N__3197),
            .I(\seq.counter.T_RNI0T6TZ0Z_4_cascade_ ));
    CascadeMux I__379 (
            .O(N__3194),
            .I(N__3191));
    InMux I__378 (
            .O(N__3191),
            .I(N__3188));
    LocalMux I__377 (
            .O(N__3188),
            .I(N__3185));
    Span4Mux_s1_h I__376 (
            .O(N__3185),
            .I(N__3177));
    InMux I__375 (
            .O(N__3184),
            .I(N__3172));
    InMux I__374 (
            .O(N__3183),
            .I(N__3172));
    InMux I__373 (
            .O(N__3182),
            .I(N__3167));
    InMux I__372 (
            .O(N__3181),
            .I(N__3167));
    InMux I__371 (
            .O(N__3180),
            .I(N__3164));
    Odrv4 I__370 (
            .O(N__3177),
            .I(ir_out_7_rep1));
    LocalMux I__369 (
            .O(N__3172),
            .I(ir_out_7_rep1));
    LocalMux I__368 (
            .O(N__3167),
            .I(ir_out_7_rep1));
    LocalMux I__367 (
            .O(N__3164),
            .I(ir_out_7_rep1));
    InMux I__366 (
            .O(N__3155),
            .I(N__3148));
    InMux I__365 (
            .O(N__3154),
            .I(N__3145));
    InMux I__364 (
            .O(N__3153),
            .I(N__3140));
    InMux I__363 (
            .O(N__3152),
            .I(N__3140));
    InMux I__362 (
            .O(N__3151),
            .I(N__3137));
    LocalMux I__361 (
            .O(N__3148),
            .I(N__3132));
    LocalMux I__360 (
            .O(N__3145),
            .I(N__3132));
    LocalMux I__359 (
            .O(N__3140),
            .I(N__3127));
    LocalMux I__358 (
            .O(N__3137),
            .I(N__3127));
    Span4Mux_v I__357 (
            .O(N__3132),
            .I(N__3124));
    Odrv12 I__356 (
            .O(N__3127),
            .I(seq_T_2_rep1));
    Odrv4 I__355 (
            .O(N__3124),
            .I(seq_T_2_rep1));
    CascadeMux I__354 (
            .O(N__3119),
            .I(\seq.D_1_0_x_cascade_ ));
    CascadeMux I__353 (
            .O(N__3116),
            .I(ROM_OE_cascade_));
    InMux I__352 (
            .O(N__3113),
            .I(N__3110));
    LocalMux I__351 (
            .O(N__3110),
            .I(\pc.program_counter_m_2 ));
    InMux I__350 (
            .O(N__3107),
            .I(N__3103));
    InMux I__349 (
            .O(N__3106),
            .I(N__3100));
    LocalMux I__348 (
            .O(N__3103),
            .I(N__3097));
    LocalMux I__347 (
            .O(N__3100),
            .I(\pc.out_1_0_iv_0 ));
    Odrv12 I__346 (
            .O(N__3097),
            .I(\pc.out_1_0_iv_0 ));
    CascadeMux I__345 (
            .O(N__3092),
            .I(\pc.G_10_0_a11_2_1_cascade_ ));
    InMux I__344 (
            .O(N__3089),
            .I(N__3086));
    LocalMux I__343 (
            .O(N__3086),
            .I(N__3083));
    Odrv4 I__342 (
            .O(N__3083),
            .I(\pc.N_23 ));
    CascadeMux I__341 (
            .O(N__3080),
            .I(\pc.program_counter_RNO_6Z0Z_2_cascade_ ));
    InMux I__340 (
            .O(N__3077),
            .I(N__3074));
    LocalMux I__339 (
            .O(N__3074),
            .I(\pc.G_10_0_a11_5_2 ));
    CascadeMux I__338 (
            .O(N__3071),
            .I(\seq.S1_1Z0Z_0_cascade_ ));
    CascadeMux I__337 (
            .O(N__3068),
            .I(seq_S1_0_cascade_));
    InMux I__336 (
            .O(N__3065),
            .I(N__3062));
    LocalMux I__335 (
            .O(N__3062),
            .I(N__3059));
    Odrv4 I__334 (
            .O(N__3059),
            .I(\pc.N_16 ));
    CascadeMux I__333 (
            .O(N__3056),
            .I(\ALU_main.N_48_cascade_ ));
    CascadeMux I__332 (
            .O(N__3053),
            .I(alu_out_m_7_cascade_));
    CascadeMux I__331 (
            .O(N__3050),
            .I(acc_out_m_7_cascade_));
    IoInMux I__330 (
            .O(N__3047),
            .I(N__3044));
    LocalMux I__329 (
            .O(N__3044),
            .I(N__3041));
    Span12Mux_s1_h I__328 (
            .O(N__3041),
            .I(N__3038));
    Odrv12 I__327 (
            .O(N__3038),
            .I(out_c_7));
    InMux I__326 (
            .O(N__3035),
            .I(N__3032));
    LocalMux I__325 (
            .O(N__3032),
            .I(\pc.out_1_2_iv_0 ));
    CascadeMux I__324 (
            .O(N__3029),
            .I(\pc.program_counter_RNO_7Z0Z_0_cascade_ ));
    InMux I__323 (
            .O(N__3026),
            .I(N__3023));
    LocalMux I__322 (
            .O(N__3023),
            .I(\pc.program_counter_RNO_3Z0Z_0 ));
    InMux I__321 (
            .O(N__3020),
            .I(N__3017));
    LocalMux I__320 (
            .O(N__3017),
            .I(\pc.program_counter_RNO_8Z0Z_0 ));
    CascadeMux I__319 (
            .O(N__3014),
            .I(\pc.program_counter_m_0_2_cascade_ ));
    CascadeMux I__318 (
            .O(N__3011),
            .I(N__3008));
    InMux I__317 (
            .O(N__3008),
            .I(N__3002));
    InMux I__316 (
            .O(N__3007),
            .I(N__3002));
    LocalMux I__315 (
            .O(N__3002),
            .I(AR_out_2));
    CascadeMux I__314 (
            .O(N__2999),
            .I(N__2995));
    InMux I__313 (
            .O(N__2998),
            .I(N__2992));
    InMux I__312 (
            .O(N__2995),
            .I(N__2989));
    LocalMux I__311 (
            .O(N__2992),
            .I(AR_out_0));
    LocalMux I__310 (
            .O(N__2989),
            .I(AR_out_0));
    InMux I__309 (
            .O(N__2984),
            .I(N__2981));
    LocalMux I__308 (
            .O(N__2981),
            .I(mem_data_2_7_0__N_7_0));
    InMux I__307 (
            .O(N__2978),
            .I(N__2975));
    LocalMux I__306 (
            .O(N__2975),
            .I(\pc.program_counter_m_0_0 ));
    CascadeMux I__305 (
            .O(N__2972),
            .I(\pc.out_1_2_iv_0_cascade_ ));
    CascadeMux I__304 (
            .O(N__2969),
            .I(\pc.tbuf.g0Z0Z_1_cascade_ ));
    InMux I__303 (
            .O(N__2966),
            .I(N__2963));
    LocalMux I__302 (
            .O(N__2963),
            .I(bus_0));
    InMux I__301 (
            .O(N__2960),
            .I(N__2957));
    LocalMux I__300 (
            .O(N__2957),
            .I(mem_data_2_7_0__N_14_0));
    CascadeMux I__299 (
            .O(N__2954),
            .I(bus_6_cascade_));
    CascadeMux I__298 (
            .O(N__2951),
            .I(N_5_0_cascade_));
    InMux I__297 (
            .O(N__2948),
            .I(N__2945));
    LocalMux I__296 (
            .O(N__2945),
            .I(N__2942));
    Span4Mux_v I__295 (
            .O(N__2942),
            .I(N__2939));
    Odrv4 I__294 (
            .O(N__2939),
            .I(mem_data_2_7_0__g1));
    CascadeMux I__293 (
            .O(N__2936),
            .I(seq_un1_IR_OE_4_1_cascade_));
    InMux I__292 (
            .O(N__2933),
            .I(N__2930));
    LocalMux I__291 (
            .O(N__2930),
            .I(N__2927));
    Span4Mux_h I__290 (
            .O(N__2927),
            .I(N__2924));
    Odrv4 I__289 (
            .O(N__2924),
            .I(\pc.program_counter_RNO_5Z0Z_0 ));
    CascadeMux I__288 (
            .O(N__2921),
            .I(\seq.un17_IR_OE_cascade_ ));
    CascadeMux I__287 (
            .O(N__2918),
            .I(seq_PC_LD_0_0_cascade_));
    InMux I__286 (
            .O(N__2915),
            .I(N__2912));
    LocalMux I__285 (
            .O(N__2912),
            .I(\seq.D_6_x ));
    CascadeMux I__284 (
            .O(N__2909),
            .I(\pc.program_counter_m_3_cascade_ ));
    InMux I__283 (
            .O(N__2906),
            .I(N__2903));
    LocalMux I__282 (
            .O(N__2903),
            .I(\pc.tbuf.gZ0Z3 ));
    CascadeMux I__281 (
            .O(N__2900),
            .I(\pc.tbuf.g0Z0Z_3_cascade_ ));
    CascadeMux I__280 (
            .O(N__2897),
            .I(bus_3_cascade_));
    CascadeMux I__279 (
            .O(N__2894),
            .I(N__2891));
    InMux I__278 (
            .O(N__2891),
            .I(N__2888));
    LocalMux I__277 (
            .O(N__2888),
            .I(N__2885));
    Odrv4 I__276 (
            .O(N__2885),
            .I(seq_MAR_LD_1_0));
    CascadeMux I__275 (
            .O(N__2882),
            .I(N__2879));
    InMux I__274 (
            .O(N__2879),
            .I(N__2876));
    LocalMux I__273 (
            .O(N__2876),
            .I(\pc.program_counter_m_3 ));
    CascadeMux I__272 (
            .O(N__2873),
            .I(\seq.DZ0Z_0_cascade_ ));
    InMux I__271 (
            .O(N__2870),
            .I(N__2867));
    LocalMux I__270 (
            .O(N__2867),
            .I(clk_c));
    IoInMux I__269 (
            .O(N__2864),
            .I(N__2861));
    LocalMux I__268 (
            .O(N__2861),
            .I(buf_clk_1));
    CascadeMux I__267 (
            .O(N__2858),
            .I(\pc.N_21_0_cascade_ ));
    CascadeMux I__266 (
            .O(N__2855),
            .I(seq_D_6_cascade_));
    InMux I__265 (
            .O(N__2852),
            .I(N__2849));
    LocalMux I__264 (
            .O(N__2849),
            .I(\pc.G_12_i_a3_1 ));
    INV \INVout_reg.ff4.qC  (
            .O(\INVout_reg.ff4.qC_net ),
            .I(N__4804));
    INV \INVb_reg.ff4.qC  (
            .O(\INVb_reg.ff4.qC_net ),
            .I(N__4807));
    INV \INVout_reg.ff2.qC  (
            .O(\INVout_reg.ff2.qC_net ),
            .I(N__4803));
    INV \INVb_reg.ff3.qC  (
            .O(\INVb_reg.ff3.qC_net ),
            .I(N__4799));
    INV \INVIR.ff1.q_nerC  (
            .O(\INVIR.ff1.q_nerC_net ),
            .I(N__4795));
    INV \INVout_reg.ff3.qC  (
            .O(\INVout_reg.ff3.qC_net ),
            .I(N__4788));
    INV \INVout_reg.ff6.qC  (
            .O(\INVout_reg.ff6.qC_net ),
            .I(N__4808));
    INV \INVb_reg.ff2.qC  (
            .O(\INVb_reg.ff2.qC_net ),
            .I(N__4806));
    INV \INVout_reg.ff7.qC  (
            .O(\INVout_reg.ff7.qC_net ),
            .I(N__4802));
    INV \INVb_reg.ff6.qC  (
            .O(\INVb_reg.ff6.qC_net ),
            .I(N__4798));
    INV \INVmar.ff4.q_nerC  (
            .O(\INVmar.ff4.q_nerC_net ),
            .I(N__4794));
    INV \INVacc.ff1.qC  (
            .O(\INVacc.ff1.qC_net ),
            .I(N__4791));
    INV \INVIR.ff2.q_nerC  (
            .O(\INVIR.ff2.q_nerC_net ),
            .I(N__4783));
    INV \INVacc.ff7.qC  (
            .O(\INVacc.ff7.qC_net ),
            .I(N__4801));
    INV \INVb_reg.ff5.qC  (
            .O(\INVb_reg.ff5.qC_net ),
            .I(N__4797));
    INV \INVAR.ff2.qC  (
            .O(\INVAR.ff2.qC_net ),
            .I(N__4779));
    INV \INVseq.q_retC  (
            .O(\INVseq.q_retC_net ),
            .I(N__4805));
    INV \INVseq.q_ret_1C  (
            .O(\INVseq.q_ret_1C_net ),
            .I(N__4800));
    INV \INVseq.counter.T_0C  (
            .O(\INVseq.counter.T_0C_net ),
            .I(N__4782));
    INV \INVIR.ff7.q_0_nerC  (
            .O(\INVIR.ff7.q_0_nerC_net ),
            .I(N__4793));
    INV \INVseq.counter.T_0_fast_2C  (
            .O(\INVseq.counter.T_0_fast_2C_net ),
            .I(N__4790));
    INV \INVIR.ff6.q_ret_1C  (
            .O(\INVIR.ff6.q_ret_1C_net ),
            .I(N__4785));
    INV \INVIR.ff7.q_0_fastC  (
            .O(\INVIR.ff7.q_0_fastC_net ),
            .I(N__4781));
    INV \INVmar.ff1.q_nerC  (
            .O(\INVmar.ff1.q_nerC_net ),
            .I(N__4778));
    INV \INVout_reg.ff8.qC  (
            .O(\INVout_reg.ff8.qC_net ),
            .I(N__4776));
    INV \INVAR.ff3.qC  (
            .O(\INVAR.ff3.qC_net ),
            .I(N__4777));
    INV \INVseq.counter.T_4C  (
            .O(\INVseq.counter.T_4C_net ),
            .I(N__4792));
    INV \INVIR.ff5.q_0_nerC  (
            .O(\INVIR.ff5.q_0_nerC_net ),
            .I(N__4789));
    INV \INVIR.ff7.q_ret_1C  (
            .O(\INVIR.ff7.q_ret_1C_net ),
            .I(N__4784));
    INV \INVIR.ff5.q_0_rep1C  (
            .O(\INVIR.ff5.q_0_rep1C_net ),
            .I(N__4780));
    INV \INVAR.ff4.qC  (
            .O(\INVAR.ff4.qC_net ),
            .I(N__4775));
    INV \INVseq.counter.T_0_2_rep1C  (
            .O(\INVseq.counter.T_0_2_rep1C_net ),
            .I(N__4774));
    defparam IN_MUX_bfv_4_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_12_0_));
    defparam IN_MUX_bfv_4_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_13_0_ (
            .carryinitin(\ALU_main.un1_A_cry_6 ),
            .carryinitout(bfn_4_13_0_));
    ICE_GB buf_clk_1_inferred_clock_0_RNIEA29 (
            .USERSIGNALTOGLOBALBUFFER(N__2864),
            .GLOBALBUFFEROUTPUT(buf_clk_1_g));
    GND GND (
            .Y(GNDG0));
    VCC VCC (
            .Y(VCCG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam \seq.counter.T_0_2_rep1_LC_1_8_0 .C_ON=1'b0;
    defparam \seq.counter.T_0_2_rep1_LC_1_8_0 .SEQ_MODE=4'b1010;
    defparam \seq.counter.T_0_2_rep1_LC_1_8_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \seq.counter.T_0_2_rep1_LC_1_8_0  (
            .in0(N__8666),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(seq_T_2_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVseq.counter.T_0_2_rep1C_net ),
            .ce(),
            .sr(N__7288));
    defparam \AR.ff1.q_LC_1_8_6 .C_ON=1'b0;
    defparam \AR.ff1.q_LC_1_8_6 .SEQ_MODE=4'b1010;
    defparam \AR.ff1.q_LC_1_8_6 .LUT_INIT=16'b1110110001001100;
    LogicCell40 \AR.ff1.q_LC_1_8_6  (
            .in0(N__4273),
            .in1(N__2998),
            .in2(N__4668),
            .in3(N__2966),
            .lcout(AR_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVseq.counter.T_0_2_rep1C_net ),
            .ce(),
            .sr(N__7288));
    defparam \seq.counter.T_0_2_LC_1_8_7 .C_ON=1'b0;
    defparam \seq.counter.T_0_2_LC_1_8_7 .SEQ_MODE=4'b1010;
    defparam \seq.counter.T_0_2_LC_1_8_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \seq.counter.T_0_2_LC_1_8_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8665),
            .lcout(seq_T_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVseq.counter.T_0_2_rep1C_net ),
            .ce(),
            .sr(N__7288));
    defparam buf_clk_1_inferred_clock_0_RNO_LC_1_9_0.C_ON=1'b0;
    defparam buf_clk_1_inferred_clock_0_RNO_LC_1_9_0.SEQ_MODE=4'b0000;
    defparam buf_clk_1_inferred_clock_0_RNO_LC_1_9_0.LUT_INIT=16'b0101010100000000;
    LogicCell40 buf_clk_1_inferred_clock_0_RNO_LC_1_9_0 (
            .in0(N__4337),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2870),
            .lcout(buf_clk_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNI1BHH1_0_LC_1_9_1 .C_ON=1'b0;
    defparam \pc.program_counter_RNI1BHH1_0_LC_1_9_1 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNI1BHH1_0_LC_1_9_1 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \pc.program_counter_RNI1BHH1_0_LC_1_9_1  (
            .in0(N__3643),
            .in1(N__4639),
            .in2(N__3548),
            .in3(N__4252),
            .lcout(\pc.program_counter_m_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_4_0_LC_1_9_3 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_4_0_LC_1_9_3 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_4_0_LC_1_9_3 .LUT_INIT=16'b0001010100000000;
    LogicCell40 \pc.program_counter_RNO_4_0_LC_1_9_3  (
            .in0(N__3541),
            .in1(N__4251),
            .in2(N__4654),
            .in3(N__4205),
            .lcout(),
            .ltout(\pc.N_21_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_1_0_LC_1_9_4 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_1_0_LC_1_9_4 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_1_0_LC_1_9_4 .LUT_INIT=16'b0101000100000000;
    LogicCell40 \pc.program_counter_RNO_1_0_LC_1_9_4  (
            .in0(N__8672),
            .in1(N__3644),
            .in2(N__2858),
            .in3(N__2933),
            .lcout(\pc.G_12_i_a3_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \mar.ff1.q_sbtinv_LC_1_9_7 .C_ON=1'b0;
    defparam \mar.ff1.q_sbtinv_LC_1_9_7 .SEQ_MODE=4'b0000;
    defparam \mar.ff1.q_sbtinv_LC_1_9_7 .LUT_INIT=16'b1010111011111111;
    LogicCell40 \mar.ff1.q_sbtinv_LC_1_9_7  (
            .in0(N__3545),
            .in1(N__4640),
            .in2(N__2894),
            .in3(N__4497),
            .lcout(\mar.MAR_LD_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_10_2_LC_1_10_0 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_10_2_LC_1_10_0 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_10_2_LC_1_10_0 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \pc.program_counter_RNO_10_2_LC_1_10_0  (
            .in0(N__3718),
            .in1(N__3152),
            .in2(N__3537),
            .in3(N__4248),
            .lcout(\pc.program_counter_m_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.decoder.D_6_LC_1_10_1 .C_ON=1'b0;
    defparam \seq.decoder.D_6_LC_1_10_1 .SEQ_MODE=4'b0000;
    defparam \seq.decoder.D_6_LC_1_10_1 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \seq.decoder.D_6_LC_1_10_1  (
            .in0(N__5455),
            .in1(N__3302),
            .in2(N__3194),
            .in3(N__5408),
            .lcout(seq_D_6),
            .ltout(seq_D_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNI0GCL1_1_LC_1_10_2 .C_ON=1'b0;
    defparam \pc.program_counter_RNI0GCL1_1_LC_1_10_2 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNI0GCL1_1_LC_1_10_2 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \pc.program_counter_RNI0GCL1_1_LC_1_10_2  (
            .in0(N__3523),
            .in1(N__4837),
            .in2(N__2855),
            .in3(N__3153),
            .lcout(\pc.program_counter_m_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_0_LC_1_10_5 .C_ON=1'b0;
    defparam \pc.program_counter_0_LC_1_10_5 .SEQ_MODE=4'b1010;
    defparam \pc.program_counter_0_LC_1_10_5 .LUT_INIT=16'b0000000101010101;
    LogicCell40 \pc.program_counter_0_LC_1_10_5  (
            .in0(N__3239),
            .in1(N__2852),
            .in2(N__3590),
            .in3(N__3026),
            .lcout(\pc.program_counterZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4773),
            .ce(),
            .sr(N__7287));
    defparam \pc.tbuf.g3_LC_1_11_1 .C_ON=1'b0;
    defparam \pc.tbuf.g3_LC_1_11_1 .SEQ_MODE=4'b0000;
    defparam \pc.tbuf.g3_LC_1_11_1 .LUT_INIT=16'b0000000001110111;
    LogicCell40 \pc.tbuf.g3_LC_1_11_1  (
            .in0(N__2948),
            .in1(N__7121),
            .in2(_gnd_net_),
            .in3(N__6482),
            .lcout(\pc.tbuf.gZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNI2ICL1_3_LC_1_11_2 .C_ON=1'b0;
    defparam \pc.program_counter_RNI2ICL1_3_LC_1_11_2 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNI2ICL1_3_LC_1_11_2 .LUT_INIT=16'b1010100010100000;
    LogicCell40 \pc.program_counter_RNI2ICL1_3_LC_1_11_2  (
            .in0(N__4009),
            .in1(N__4249),
            .in2(N__3547),
            .in3(N__3155),
            .lcout(\pc.program_counter_m_3 ),
            .ltout(\pc.program_counter_m_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.tbuf.g0_3_LC_1_11_3 .C_ON=1'b0;
    defparam \pc.tbuf.g0_3_LC_1_11_3 .SEQ_MODE=4'b0000;
    defparam \pc.tbuf.g0_3_LC_1_11_3 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \pc.tbuf.g0_3_LC_1_11_3  (
            .in0(N__4485),
            .in1(N__3890),
            .in2(N__2909),
            .in3(N__2906),
            .lcout(\pc.tbuf.g0Z0Z_3 ),
            .ltout(\pc.tbuf.g0Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.tbuf.g0_LC_1_11_4 .C_ON=1'b0;
    defparam \pc.tbuf.g0_LC_1_11_4 .SEQ_MODE=4'b0000;
    defparam \pc.tbuf.g0_LC_1_11_4 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \pc.tbuf.g0_LC_1_11_4  (
            .in0(N__7618),
            .in1(N__7749),
            .in2(N__2900),
            .in3(N__7544),
            .lcout(),
            .ltout(bus_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \AR.ff4.q_LC_1_11_5 .C_ON=1'b0;
    defparam \AR.ff4.q_LC_1_11_5 .SEQ_MODE=4'b1010;
    defparam \AR.ff4.q_LC_1_11_5 .LUT_INIT=16'b1110010011001100;
    LogicCell40 \AR.ff4.q_LC_1_11_5  (
            .in0(N__4250),
            .in1(N__3912),
            .in2(N__2897),
            .in3(N__4669),
            .lcout(\AR.ff4.AR_out_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVAR.ff4.qC_net ),
            .ce(),
            .sr(N__7289));
    defparam \seq.MAR_LD_1_0_LC_1_12_0 .C_ON=1'b0;
    defparam \seq.MAR_LD_1_0_LC_1_12_0 .SEQ_MODE=4'b0000;
    defparam \seq.MAR_LD_1_0_LC_1_12_0 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \seq.MAR_LD_1_0_LC_1_12_0  (
            .in0(N__4965),
            .in1(N__5138),
            .in2(_gnd_net_),
            .in3(N__5005),
            .lcout(seq_MAR_LD_1_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.g2_0_LC_1_12_1 .C_ON=1'b0;
    defparam \seq.g2_0_LC_1_12_1 .SEQ_MODE=4'b0000;
    defparam \seq.g2_0_LC_1_12_1 .LUT_INIT=16'b0000000000000101;
    LogicCell40 \seq.g2_0_LC_1_12_1  (
            .in0(N__5004),
            .in1(_gnd_net_),
            .in2(N__5147),
            .in3(N__4964),
            .lcout(\seq.g2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.tbuf.out_1_iv_1_1_LC_1_12_2 .C_ON=1'b0;
    defparam \pc.tbuf.out_1_iv_1_1_LC_1_12_2 .SEQ_MODE=4'b0000;
    defparam \pc.tbuf.out_1_iv_1_1_LC_1_12_2 .LUT_INIT=16'b0000101100000011;
    LogicCell40 \pc.tbuf.out_1_iv_1_1_LC_1_12_2  (
            .in0(N__3328),
            .in1(N__3888),
            .in2(N__2882),
            .in3(N__4541),
            .lcout(\pc.out_1_iv_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.decoder.D_0_LC_1_12_3 .C_ON=1'b0;
    defparam \seq.decoder.D_0_LC_1_12_3 .SEQ_MODE=4'b0000;
    defparam \seq.decoder.D_0_LC_1_12_3 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \seq.decoder.D_0_LC_1_12_3  (
            .in0(N__3434),
            .in1(N__3272),
            .in2(N__3215),
            .in3(N__5500),
            .lcout(\seq.DZ0Z_0 ),
            .ltout(\seq.DZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_0_2_rep1_RNIE27K3_LC_1_12_4 .C_ON=1'b0;
    defparam \seq.counter.T_0_2_rep1_RNIE27K3_LC_1_12_4 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_0_2_rep1_RNIE27K3_LC_1_12_4 .LUT_INIT=16'b0101010101010111;
    LogicCell40 \seq.counter.T_0_2_rep1_RNIE27K3_LC_1_12_4  (
            .in0(N__3151),
            .in1(N__5134),
            .in2(N__2873),
            .in3(N__5003),
            .lcout(seq_un1_IR_OE_4_1),
            .ltout(seq_un1_IR_OE_4_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_3_2_LC_1_12_5 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_3_2_LC_1_12_5 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_3_2_LC_1_12_5 .LUT_INIT=16'b0111111101010101;
    LogicCell40 \pc.program_counter_RNO_3_2_LC_1_12_5  (
            .in0(N__4539),
            .in1(N__4457),
            .in2(N__2936),
            .in3(N__4194),
            .lcout(\pc.G_10_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_5_0_LC_1_12_7 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_5_0_LC_1_12_7 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_5_0_LC_1_12_7 .LUT_INIT=16'b1000111100001111;
    LogicCell40 \pc.program_counter_RNO_5_0_LC_1_12_7  (
            .in0(N__4540),
            .in1(N__3327),
            .in2(N__8765),
            .in3(N__4458),
            .lcout(\pc.program_counter_RNO_5Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_8_2_LC_1_13_0 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_8_2_LC_1_13_0 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_8_2_LC_1_13_0 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \pc.program_counter_RNO_8_2_LC_1_13_0  (
            .in0(N__8667),
            .in1(N__4547),
            .in2(N__3722),
            .in3(N__4183),
            .lcout(\pc.N_23 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.q_ret_RNI7NFN_LC_1_13_1 .C_ON=1'b0;
    defparam \seq.q_ret_RNI7NFN_LC_1_13_1 .SEQ_MODE=4'b0000;
    defparam \seq.q_ret_RNI7NFN_LC_1_13_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \seq.q_ret_RNI7NFN_LC_1_13_1  (
            .in0(N__3184),
            .in1(N__5561),
            .in2(N__4292),
            .in3(N__5398),
            .lcout(),
            .ltout(\seq.un17_IR_OE_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_RNIPKHM1_3_LC_1_13_2 .C_ON=1'b0;
    defparam \seq.counter.T_RNIPKHM1_3_LC_1_13_2 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_RNIPKHM1_3_LC_1_13_2 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \seq.counter.T_RNIPKHM1_3_LC_1_13_2  (
            .in0(N__5218),
            .in1(N__2915),
            .in2(N__2921),
            .in3(N__3301),
            .lcout(seq_PC_LD_0_0),
            .ltout(seq_PC_LD_0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_0_3_LC_1_13_3 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_0_3_LC_1_13_3 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_0_3_LC_1_13_3 .LUT_INIT=16'b1100110011101111;
    LogicCell40 \pc.program_counter_RNO_0_3_LC_1_13_3  (
            .in0(N__4184),
            .in1(N__3560),
            .in2(N__2918),
            .in3(N__8668),
            .lcout(\pc.g0_rn_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.decoder.D_6_x_LC_1_13_4 .C_ON=1'b0;
    defparam \seq.decoder.D_6_x_LC_1_13_4 .SEQ_MODE=4'b0000;
    defparam \seq.decoder.D_6_x_LC_1_13_4 .LUT_INIT=16'b0000000000100010;
    LogicCell40 \seq.decoder.D_6_x_LC_1_13_4  (
            .in0(N__5397),
            .in1(N__5443),
            .in2(_gnd_net_),
            .in3(N__3183),
            .lcout(\seq.D_6_x ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \IR.ff5.q_0_rep1_LC_1_13_6 .C_ON=1'b0;
    defparam \IR.ff5.q_0_rep1_LC_1_13_6 .SEQ_MODE=4'b1010;
    defparam \IR.ff5.q_0_rep1_LC_1_13_6 .LUT_INIT=16'b1111101000001010;
    LogicCell40 \IR.ff5.q_0_rep1_LC_1_13_6  (
            .in0(N__5562),
            .in1(_gnd_net_),
            .in2(N__8686),
            .in3(N__5594),
            .lcout(ir_out_4_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVIR.ff5.q_0_rep1C_net ),
            .ce(),
            .sr(N__7294));
    defparam \seq.decoder.D_4_0_LC_1_13_7 .C_ON=1'b0;
    defparam \seq.decoder.D_4_0_LC_1_13_7 .SEQ_MODE=4'b0000;
    defparam \seq.decoder.D_4_0_LC_1_13_7 .LUT_INIT=16'b0000000001000000;
    LogicCell40 \seq.decoder.D_4_0_LC_1_13_7  (
            .in0(N__5444),
            .in1(N__5494),
            .in2(N__5407),
            .in3(N__3180),
            .lcout(\seq.D_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buf1.out_1_0_iv_LC_1_14_1 .C_ON=1'b0;
    defparam \buf1.out_1_0_iv_LC_1_14_1 .SEQ_MODE=4'b0000;
    defparam \buf1.out_1_0_iv_LC_1_14_1 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \buf1.out_1_0_iv_LC_1_14_1  (
            .in0(N__6829),
            .in1(N__6789),
            .in2(N__6746),
            .in3(N__6521),
            .lcout(bus_6),
            .ltout(bus_6_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \IR.ff7.q_0_ner_RNI7C4KI_LC_1_14_2 .C_ON=1'b0;
    defparam \IR.ff7.q_0_ner_RNI7C4KI_LC_1_14_2 .SEQ_MODE=4'b0000;
    defparam \IR.ff7.q_0_ner_RNI7C4KI_LC_1_14_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \IR.ff7.q_0_ner_RNI7C4KI_LC_1_14_2  (
            .in0(_gnd_net_),
            .in1(N__8660),
            .in2(N__2954),
            .in3(N__3964),
            .lcout(N_5_0),
            .ltout(N_5_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \IR.ff7.q_ret_1_LC_1_14_3 .C_ON=1'b0;
    defparam \IR.ff7.q_ret_1_LC_1_14_3 .SEQ_MODE=4'b1011;
    defparam \IR.ff7.q_ret_1_LC_1_14_3 .LUT_INIT=16'b0000111100001111;
    LogicCell40 \IR.ff7.q_ret_1_LC_1_14_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2951),
            .in3(_gnd_net_),
            .lcout(ir_out_i_2_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVIR.ff7.q_ret_1C_net ),
            .ce(),
            .sr(N__7298));
    defparam \seq.g0_i_a3_2_LC_1_14_4 .C_ON=1'b0;
    defparam \seq.g0_i_a3_2_LC_1_14_4 .SEQ_MODE=4'b0000;
    defparam \seq.g0_i_a3_2_LC_1_14_4 .LUT_INIT=16'b0100010000000000;
    LogicCell40 \seq.g0_i_a3_2_LC_1_14_4  (
            .in0(N__5545),
            .in1(N__3295),
            .in2(_gnd_net_),
            .in3(N__3374),
            .lcout(\seq.g0_i_a3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \IR.ff6.q_0_fast_LC_1_14_5 .C_ON=1'b0;
    defparam \IR.ff6.q_0_fast_LC_1_14_5 .SEQ_MODE=4'b1010;
    defparam \IR.ff6.q_0_fast_LC_1_14_5 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \IR.ff6.q_0_fast_LC_1_14_5  (
            .in0(N__8661),
            .in1(N__6086),
            .in2(_gnd_net_),
            .in3(N__4417),
            .lcout(IR_ff6_q_0_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVIR.ff7.q_ret_1C_net ),
            .ce(),
            .sr(N__7298));
    defparam \seq.decoder.D_3_0_LC_1_14_6 .C_ON=1'b0;
    defparam \seq.decoder.D_3_0_LC_1_14_6 .SEQ_MODE=4'b0000;
    defparam \seq.decoder.D_3_0_LC_1_14_6 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \seq.decoder.D_3_0_LC_1_14_6  (
            .in0(N__5445),
            .in1(N__3296),
            .in2(N__3424),
            .in3(N__3265),
            .lcout(\seq.D_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \IR.ff7.q_ret_1_fast_LC_1_14_7 .C_ON=1'b0;
    defparam \IR.ff7.q_ret_1_fast_LC_1_14_7 .SEQ_MODE=4'b1011;
    defparam \IR.ff7.q_ret_1_fast_LC_1_14_7 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \IR.ff7.q_ret_1_fast_LC_1_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4351),
            .lcout(IR_ff7_q_ret_1_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVIR.ff7.q_ret_1C_net ),
            .ce(),
            .sr(N__7298));
    defparam \IR.ff5.q_0_ner_LC_1_15_5 .C_ON=1'b0;
    defparam \IR.ff5.q_0_ner_LC_1_15_5 .SEQ_MODE=4'b1010;
    defparam \IR.ff5.q_0_ner_LC_1_15_5 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \IR.ff5.q_0_ner_LC_1_15_5  (
            .in0(N__7995),
            .in1(N__7964),
            .in2(N__7922),
            .in3(N__7388),
            .lcout(ir_out_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVIR.ff5.q_0_nerC_net ),
            .ce(N__8683),
            .sr(N__7303));
    defparam \seq.counter.T_4_LC_1_16_0 .C_ON=1'b0;
    defparam \seq.counter.T_4_LC_1_16_0 .SEQ_MODE=4'b1010;
    defparam \seq.counter.T_4_LC_1_16_0 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \seq.counter.T_4_LC_1_16_0  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5222),
            .lcout(\seq.counter.TZ0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVseq.counter.T_4C_net ),
            .ce(),
            .sr(N__7306));
    defparam \mem.data_2_7_0__g1_LC_2_7_7 .C_ON=1'b0;
    defparam \mem.data_2_7_0__g1_LC_2_7_7 .SEQ_MODE=4'b0000;
    defparam \mem.data_2_7_0__g1_LC_2_7_7 .LUT_INIT=16'b0110011011101110;
    LogicCell40 \mem.data_2_7_0__g1_LC_2_7_7  (
            .in0(N__7044),
            .in1(N__7186),
            .in2(_gnd_net_),
            .in3(N__6965),
            .lcout(mem_data_2_7_0__g1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.tbuf.out_1_0_iv_0_LC_2_8_0 .C_ON=1'b0;
    defparam \pc.tbuf.out_1_0_iv_0_LC_2_8_0 .SEQ_MODE=4'b0000;
    defparam \pc.tbuf.out_1_0_iv_0_LC_2_8_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \pc.tbuf.out_1_0_iv_0_LC_2_8_0  (
            .in0(N__3007),
            .in1(N__4204),
            .in2(N__5993),
            .in3(N__7441),
            .lcout(\pc.out_1_0_iv_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNI3DHH1_2_LC_2_8_1 .C_ON=1'b0;
    defparam \pc.program_counter_RNI3DHH1_2_LC_2_8_1 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNI3DHH1_2_LC_2_8_1 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \pc.program_counter_RNI3DHH1_2_LC_2_8_1  (
            .in0(N__3546),
            .in1(N__3711),
            .in2(N__4666),
            .in3(N__4271),
            .lcout(),
            .ltout(\pc.program_counter_m_0_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.tbuf.g0_9_LC_2_8_2 .C_ON=1'b0;
    defparam \pc.tbuf.g0_9_LC_2_8_2 .SEQ_MODE=4'b0000;
    defparam \pc.tbuf.g0_9_LC_2_8_2 .LUT_INIT=16'b1111110011111101;
    LogicCell40 \pc.tbuf.g0_9_LC_2_8_2  (
            .in0(N__2960),
            .in1(N__3106),
            .in2(N__3014),
            .in3(N__6522),
            .lcout(\pc.tbuf.g0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \AR.ff3.q_LC_2_8_4 .C_ON=1'b0;
    defparam \AR.ff3.q_LC_2_8_4 .SEQ_MODE=4'b1010;
    defparam \AR.ff3.q_LC_2_8_4 .LUT_INIT=16'b1111100001110000;
    LogicCell40 \AR.ff3.q_LC_2_8_4  (
            .in0(N__4272),
            .in1(N__4644),
            .in2(N__3011),
            .in3(N__3455),
            .lcout(AR_out_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVAR.ff3.qC_net ),
            .ce(),
            .sr(N__7291));
    defparam \mem.data_2_7_0__g0_2_LC_2_9_0 .C_ON=1'b0;
    defparam \mem.data_2_7_0__g0_2_LC_2_9_0 .SEQ_MODE=4'b0000;
    defparam \mem.data_2_7_0__g0_2_LC_2_9_0 .LUT_INIT=16'b0111111110110101;
    LogicCell40 \mem.data_2_7_0__g0_2_LC_2_9_0  (
            .in0(N__7130),
            .in1(N__7057),
            .in2(N__7196),
            .in3(N__6967),
            .lcout(mem_data_2_7_0__N_7_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.tbuf.out_1_2_iv_0_LC_2_9_1 .C_ON=1'b0;
    defparam \pc.tbuf.out_1_2_iv_0_LC_2_9_1 .SEQ_MODE=4'b0000;
    defparam \pc.tbuf.out_1_2_iv_0_LC_2_9_1 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \pc.tbuf.out_1_2_iv_0_LC_2_9_1  (
            .in0(N__6067),
            .in1(N__4203),
            .in2(N__2999),
            .in3(N__7398),
            .lcout(\pc.out_1_2_iv_0 ),
            .ltout(\pc.out_1_2_iv_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.tbuf.g0_5_LC_2_9_2 .C_ON=1'b0;
    defparam \pc.tbuf.g0_5_LC_2_9_2 .SEQ_MODE=4'b0000;
    defparam \pc.tbuf.g0_5_LC_2_9_2 .LUT_INIT=16'b1111110011111101;
    LogicCell40 \pc.tbuf.g0_5_LC_2_9_2  (
            .in0(N__2984),
            .in1(N__2978),
            .in2(N__2972),
            .in3(N__6523),
            .lcout(\pc.tbuf.g0Z0Z_1 ),
            .ltout(\pc.tbuf.g0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.tbuf.g0_4_LC_2_9_3 .C_ON=1'b0;
    defparam \pc.tbuf.g0_4_LC_2_9_3 .SEQ_MODE=4'b0000;
    defparam \pc.tbuf.g0_4_LC_2_9_3 .LUT_INIT=16'b1111111111110100;
    LogicCell40 \pc.tbuf.g0_4_LC_2_9_3  (
            .in0(N__8877),
            .in1(N__8764),
            .in2(N__2969),
            .in3(N__8814),
            .lcout(bus_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \mem.data_2_7_0__g0_3_LC_2_9_7 .C_ON=1'b0;
    defparam \mem.data_2_7_0__g0_3_LC_2_9_7 .SEQ_MODE=4'b0000;
    defparam \mem.data_2_7_0__g0_3_LC_2_9_7 .LUT_INIT=16'b0111111110100111;
    LogicCell40 \mem.data_2_7_0__g0_3_LC_2_9_7  (
            .in0(N__6966),
            .in1(N__7192),
            .in2(N__7058),
            .in3(N__7129),
            .lcout(mem_data_2_7_0__N_14_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.ALU_Out_0_7_LC_2_10_0 .C_ON=1'b0;
    defparam \ALU_main.ALU_Out_0_7_LC_2_10_0 .SEQ_MODE=4'b0000;
    defparam \ALU_main.ALU_Out_0_7_LC_2_10_0 .LUT_INIT=16'b1000100001100110;
    LogicCell40 \ALU_main.ALU_Out_0_7_LC_2_10_0  (
            .in0(N__6269),
            .in1(N__5875),
            .in2(_gnd_net_),
            .in3(N__6194),
            .lcout(),
            .ltout(\ALU_main.N_48_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.un1_A_cry_6_c_RNIGN9C9_LC_2_10_1 .C_ON=1'b0;
    defparam \ALU_main.un1_A_cry_6_c_RNIGN9C9_LC_2_10_1 .SEQ_MODE=4'b0000;
    defparam \ALU_main.un1_A_cry_6_c_RNIGN9C9_LC_2_10_1 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \ALU_main.un1_A_cry_6_c_RNIGN9C9_LC_2_10_1  (
            .in0(N__3791),
            .in1(N__5742),
            .in2(N__3056),
            .in3(N__5644),
            .lcout(alu_out_m_7),
            .ltout(alu_out_m_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buf1.out_1_iv_LC_2_10_2 .C_ON=1'b0;
    defparam \buf1.out_1_iv_LC_2_10_2 .SEQ_MODE=4'b0000;
    defparam \buf1.out_1_iv_LC_2_10_2 .LUT_INIT=16'b1111111111110001;
    LogicCell40 \buf1.out_1_iv_LC_2_10_2  (
            .in0(N__6465),
            .in1(N__6901),
            .in2(N__3053),
            .in3(N__6327),
            .lcout(bus_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \acc.ff8.q_RNI449H1_LC_2_10_3 .C_ON=1'b0;
    defparam \acc.ff8.q_RNI449H1_LC_2_10_3 .SEQ_MODE=4'b0000;
    defparam \acc.ff8.q_RNI449H1_LC_2_10_3 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \acc.ff8.q_RNI449H1_LC_2_10_3  (
            .in0(N__5876),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7399),
            .lcout(acc_out_m_7),
            .ltout(acc_out_m_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \out_reg.ff8.q_LC_2_10_4 .C_ON=1'b0;
    defparam \out_reg.ff8.q_LC_2_10_4 .SEQ_MODE=4'b1010;
    defparam \out_reg.ff8.q_LC_2_10_4 .LUT_INIT=16'b1111110011111101;
    LogicCell40 \out_reg.ff8.q_LC_2_10_4  (
            .in0(N__6466),
            .in1(N__6293),
            .in2(N__3050),
            .in3(N__6902),
            .lcout(out_c_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVout_reg.ff8.qC_net ),
            .ce(N__7480),
            .sr(N__7290));
    defparam \pc.program_counter_RNO_7_0_LC_2_10_5 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_7_0_LC_2_10_5 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_7_0_LC_2_10_5 .LUT_INIT=16'b0011001100100010;
    LogicCell40 \pc.program_counter_RNO_7_0_LC_2_10_5  (
            .in0(N__6221),
            .in1(N__3035),
            .in2(_gnd_net_),
            .in3(N__6464),
            .lcout(),
            .ltout(\pc.program_counter_RNO_7Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_3_0_LC_2_10_6 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_3_0_LC_2_10_6 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_3_0_LC_2_10_6 .LUT_INIT=16'b0001000001010000;
    LogicCell40 \pc.program_counter_RNO_3_0_LC_2_10_6  (
            .in0(N__3065),
            .in1(N__3020),
            .in2(N__3029),
            .in3(N__5033),
            .lcout(\pc.program_counter_RNO_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_8_0_LC_2_10_7 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_8_0_LC_2_10_7 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_8_0_LC_2_10_7 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \pc.program_counter_RNO_8_0_LC_2_10_7  (
            .in0(_gnd_net_),
            .in1(N__5741),
            .in2(_gnd_net_),
            .in3(N__5643),
            .lcout(\pc.program_counter_RNO_8Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \mem.data_2_7_0__g0_LC_2_11_0 .C_ON=1'b0;
    defparam \mem.data_2_7_0__g0_LC_2_11_0 .SEQ_MODE=4'b0000;
    defparam \mem.data_2_7_0__g0_LC_2_11_0 .LUT_INIT=16'b0100100011001000;
    LogicCell40 \mem.data_2_7_0__g0_LC_2_11_0  (
            .in0(N__7174),
            .in1(N__7118),
            .in2(N__7043),
            .in3(N__6933),
            .lcout(mem_data_2_7_0__N_16_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \mar.ff1.q_ner_LC_2_11_1 .C_ON=1'b0;
    defparam \mar.ff1.q_ner_LC_2_11_1 .SEQ_MODE=4'b1010;
    defparam \mar.ff1.q_ner_LC_2_11_1 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \mar.ff1.q_ner_LC_2_11_1  (
            .in0(N__8908),
            .in1(N__8763),
            .in2(N__8878),
            .in3(N__8807),
            .lcout(mar_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVmar.ff1.q_nerC_net ),
            .ce(N__6382),
            .sr(N__7292));
    defparam \seq.counter.T_RNI4RN46_3_LC_2_11_2 .C_ON=1'b0;
    defparam \seq.counter.T_RNI4RN46_3_LC_2_11_2 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_RNI4RN46_3_LC_2_11_2 .LUT_INIT=16'b0000011100000000;
    LogicCell40 \seq.counter.T_RNI4RN46_3_LC_2_11_2  (
            .in0(N__5217),
            .in1(N__4963),
            .in2(N__8684),
            .in3(N__3311),
            .lcout(ROM_OE),
            .ltout(ROM_OE_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_7_2_LC_2_11_3 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_7_2_LC_2_11_3 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_7_2_LC_2_11_3 .LUT_INIT=16'b0000000000000100;
    LogicCell40 \pc.program_counter_RNO_7_2_LC_2_11_3  (
            .in0(N__6934),
            .in1(N__7018),
            .in2(N__3116),
            .in3(N__7120),
            .lcout(\pc.G_10_0_a11_5_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_9_2_LC_2_11_4 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_9_2_LC_2_11_4 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_9_2_LC_2_11_4 .LUT_INIT=16'b1000001000000000;
    LogicCell40 \pc.program_counter_RNO_9_2_LC_2_11_4  (
            .in0(N__7173),
            .in1(N__7119),
            .in2(N__7042),
            .in3(N__6932),
            .lcout(),
            .ltout(\pc.G_10_0_a11_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_6_2_LC_2_11_5 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_6_2_LC_2_11_5 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_6_2_LC_2_11_5 .LUT_INIT=16'b1110111011111110;
    LogicCell40 \pc.program_counter_RNO_6_2_LC_2_11_5  (
            .in0(N__3113),
            .in1(N__3107),
            .in2(N__3092),
            .in3(N__6463),
            .lcout(),
            .ltout(\pc.program_counter_RNO_6Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_2_2_LC_2_11_6 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_2_2_LC_2_11_6 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_2_2_LC_2_11_6 .LUT_INIT=16'b1110111011101010;
    LogicCell40 \pc.program_counter_RNO_2_2_LC_2_11_6  (
            .in0(N__3089),
            .in1(N__3769),
            .in2(N__3080),
            .in3(N__3077),
            .lcout(\pc.G_10_0_sx ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.S1_1_0_LC_2_12_0 .C_ON=1'b0;
    defparam \seq.S1_1_0_LC_2_12_0 .SEQ_MODE=4'b0000;
    defparam \seq.S1_1_0_LC_2_12_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \seq.S1_1_0_LC_2_12_0  (
            .in0(N__5499),
            .in1(N__3211),
            .in2(_gnd_net_),
            .in3(N__5405),
            .lcout(),
            .ltout(\seq.S1_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_RNIMQC72_4_LC_2_12_1 .C_ON=1'b0;
    defparam \seq.counter.T_RNIMQC72_4_LC_2_12_1 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_RNIMQC72_4_LC_2_12_1 .LUT_INIT=16'b0101010111011111;
    LogicCell40 \seq.counter.T_RNIMQC72_4_LC_2_12_1  (
            .in0(N__5350),
            .in1(N__3182),
            .in2(N__3071),
            .in3(N__4897),
            .lcout(seq_S1_0),
            .ltout(seq_S1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_9_0_LC_2_12_2 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_9_0_LC_2_12_2 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_9_0_LC_2_12_2 .LUT_INIT=16'b0000100100000010;
    LogicCell40 \pc.program_counter_RNO_9_0_LC_2_12_2  (
            .in0(N__6245),
            .in1(N__6186),
            .in2(N__3068),
            .in3(N__6068),
            .lcout(\pc.N_16 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \IR.ff7.q_0_fast_LC_2_12_3 .C_ON=1'b0;
    defparam \IR.ff7.q_0_fast_LC_2_12_3 .SEQ_MODE=4'b1010;
    defparam \IR.ff7.q_0_fast_LC_2_12_3 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \IR.ff7.q_0_fast_LC_2_12_3  (
            .in0(N__3967),
            .in1(N__3224),
            .in2(_gnd_net_),
            .in3(N__8663),
            .lcout(IR_ff7_q_0_fast),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVIR.ff7.q_0_fastC_net ),
            .ce(),
            .sr(N__7295));
    defparam \IR.ff5.q_0_fast_LC_2_12_4 .C_ON=1'b0;
    defparam \IR.ff5.q_0_fast_LC_2_12_4 .SEQ_MODE=4'b1010;
    defparam \IR.ff5.q_0_fast_LC_2_12_4 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \IR.ff5.q_0_fast_LC_2_12_4  (
            .in0(N__5590),
            .in1(N__8662),
            .in2(_gnd_net_),
            .in3(N__5564),
            .lcout(ir_out_fast_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVIR.ff7.q_0_fastC_net ),
            .ce(),
            .sr(N__7295));
    defparam \seq.counter.T_RNI0T6T_4_LC_2_12_5 .C_ON=1'b0;
    defparam \seq.counter.T_RNI0T6T_4_LC_2_12_5 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_RNI0T6T_4_LC_2_12_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \seq.counter.T_RNI0T6T_4_LC_2_12_5  (
            .in0(N__3210),
            .in1(N__3181),
            .in2(N__5362),
            .in3(N__5498),
            .lcout(),
            .ltout(\seq.counter.T_RNI0T6TZ0Z_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_RNI0TT62_4_LC_2_12_6 .C_ON=1'b0;
    defparam \seq.counter.T_RNI0TT62_4_LC_2_12_6 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_RNI0TT62_4_LC_2_12_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \seq.counter.T_RNI0TT62_4_LC_2_12_6  (
            .in0(N__3476),
            .in1(N__3966),
            .in2(N__3197),
            .in3(N__3386),
            .lcout(seq_S0_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \IR.ff8.q_0_rep1_LC_2_12_7 .C_ON=1'b0;
    defparam \IR.ff8.q_0_rep1_LC_2_12_7 .SEQ_MODE=4'b1010;
    defparam \IR.ff8.q_0_rep1_LC_2_12_7 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \IR.ff8.q_0_rep1_LC_2_12_7  (
            .in0(N__4383),
            .in1(N__8664),
            .in2(_gnd_net_),
            .in3(N__5311),
            .lcout(ir_out_7_rep1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVIR.ff7.q_0_fastC_net ),
            .ce(),
            .sr(N__7295));
    defparam \seq.decoder.D_1_0_x_LC_2_13_0 .C_ON=1'b0;
    defparam \seq.decoder.D_1_0_x_LC_2_13_0 .SEQ_MODE=4'b0000;
    defparam \seq.decoder.D_1_0_x_LC_2_13_0 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \seq.decoder.D_1_0_x_LC_2_13_0  (
            .in0(N__5497),
            .in1(N__3428),
            .in2(_gnd_net_),
            .in3(N__3268),
            .lcout(),
            .ltout(\seq.D_1_0_x_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_0_2_rep1_RNIC9OP2_LC_2_13_1 .C_ON=1'b0;
    defparam \seq.counter.T_0_2_rep1_RNIC9OP2_LC_2_13_1 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_0_2_rep1_RNIC9OP2_LC_2_13_1 .LUT_INIT=16'b0011011101110111;
    LogicCell40 \seq.counter.T_0_2_rep1_RNIC9OP2_LC_2_13_1  (
            .in0(N__4890),
            .in1(N__3154),
            .in2(N__3119),
            .in3(N__5448),
            .lcout(seq_MAR_LD_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \IR.ff6.q_ret_1_LC_2_13_3 .C_ON=1'b0;
    defparam \IR.ff6.q_ret_1_LC_2_13_3 .SEQ_MODE=4'b1011;
    defparam \IR.ff6.q_ret_1_LC_2_13_3 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \IR.ff6.q_ret_1_LC_2_13_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4316),
            .lcout(ir_out_i_2_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVIR.ff6.q_ret_1C_net ),
            .ce(),
            .sr(N__7299));
    defparam \seq.B_LD_2_tz_LC_2_13_4 .C_ON=1'b0;
    defparam \seq.B_LD_2_tz_LC_2_13_4 .SEQ_MODE=4'b0000;
    defparam \seq.B_LD_2_tz_LC_2_13_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \seq.B_LD_2_tz_LC_2_13_4  (
            .in0(_gnd_net_),
            .in1(N__4889),
            .in2(_gnd_net_),
            .in3(N__5002),
            .lcout(\seq.B_LD_0_2_tz ),
            .ltout(\seq.B_LD_0_2_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_RNIR83I4_0_3_LC_2_13_5 .C_ON=1'b0;
    defparam \seq.counter.T_RNIR83I4_0_3_LC_2_13_5 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_RNIR83I4_0_3_LC_2_13_5 .LUT_INIT=16'b0101010101110101;
    LogicCell40 \seq.counter.T_RNIR83I4_0_3_LC_2_13_5  (
            .in0(N__5216),
            .in1(N__5133),
            .in2(N__3314),
            .in3(N__5078),
            .lcout(\seq.counter.T_RNIR83I4_0Z0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.decoder.D_2_0_LC_2_13_6 .C_ON=1'b0;
    defparam \seq.decoder.D_2_0_LC_2_13_6 .SEQ_MODE=4'b0000;
    defparam \seq.decoder.D_2_0_LC_2_13_6 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \seq.decoder.D_2_0_LC_2_13_6  (
            .in0(N__5446),
            .in1(N__3267),
            .in2(N__3432),
            .in3(N__3297),
            .lcout(\seq.D_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.decoder.D_1_0_LC_2_13_7 .C_ON=1'b0;
    defparam \seq.decoder.D_1_0_LC_2_13_7 .SEQ_MODE=4'b0000;
    defparam \seq.decoder.D_1_0_LC_2_13_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \seq.decoder.D_1_0_LC_2_13_7  (
            .in0(N__3266),
            .in1(N__5496),
            .in2(N__3433),
            .in3(N__5447),
            .lcout(\seq.D_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_RNIGQT43_1_LC_2_14_0 .C_ON=1'b0;
    defparam \seq.counter.T_RNIGQT43_1_LC_2_14_0 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_RNIGQT43_1_LC_2_14_0 .LUT_INIT=16'b0011001100010001;
    LogicCell40 \seq.counter.T_RNIGQT43_1_LC_2_14_0  (
            .in0(N__4542),
            .in1(N__8654),
            .in2(_gnd_net_),
            .in3(N__4179),
            .lcout(N_30),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_0_fast_RNIP4D21_2_LC_2_14_1 .C_ON=1'b0;
    defparam \seq.counter.T_0_fast_RNIP4D21_2_LC_2_14_1 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_0_fast_RNIP4D21_2_LC_2_14_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \seq.counter.T_0_fast_RNIP4D21_2_LC_2_14_1  (
            .in0(N__3351),
            .in1(N__4413),
            .in2(N__3965),
            .in3(N__5290),
            .lcout(),
            .ltout(\seq.counter.T_0_fast_RNIP4D21Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_0_fast_RNILB791_2_LC_2_14_2 .C_ON=1'b0;
    defparam \seq.counter.T_0_fast_RNILB791_2_LC_2_14_2 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_0_fast_RNILB791_2_LC_2_14_2 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \seq.counter.T_0_fast_RNILB791_2_LC_2_14_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3245),
            .in3(N__5548),
            .lcout(T_0_fast_RNILB791_2),
            .ltout(T_0_fast_RNILB791_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_0_0_LC_2_14_3 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_0_0_LC_2_14_3 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_0_0_LC_2_14_3 .LUT_INIT=16'b1000100110001000;
    LogicCell40 \pc.program_counter_RNO_0_0_LC_2_14_3  (
            .in0(N__8655),
            .in1(N__3671),
            .in2(N__3242),
            .in3(N__4543),
            .lcout(\pc.G_12_i_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_0_fast_2_LC_2_14_4 .C_ON=1'b0;
    defparam \seq.counter.T_0_fast_2_LC_2_14_4 .SEQ_MODE=4'b1010;
    defparam \seq.counter.T_0_fast_2_LC_2_14_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \seq.counter.T_0_fast_2_LC_2_14_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8659),
            .lcout(\seq.counter.T_fast_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVseq.counter.T_0_fast_2C_net ),
            .ce(),
            .sr(N__7304));
    defparam \seq.counter.T_0_fast_RNIG89V_2_LC_2_14_5 .C_ON=1'b0;
    defparam \seq.counter.T_0_fast_RNIG89V_2_LC_2_14_5 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_0_fast_RNIG89V_2_LC_2_14_5 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \seq.counter.T_0_fast_RNIG89V_2_LC_2_14_5  (
            .in0(N__3377),
            .in1(N__3409),
            .in2(N__3355),
            .in3(N__5495),
            .lcout(),
            .ltout(\seq.counter.T_0_fast_RNIG89VZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_0_fast_RNICF361_2_LC_2_14_6 .C_ON=1'b0;
    defparam \seq.counter.T_0_fast_RNICF361_2_LC_2_14_6 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_0_fast_RNICF361_2_LC_2_14_6 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \seq.counter.T_0_fast_RNICF361_2_LC_2_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3227),
            .in3(N__5549),
            .lcout(OUT_LD),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \IR.ff8.q_0_fast_LC_2_14_7 .C_ON=1'b0;
    defparam \IR.ff8.q_0_fast_LC_2_14_7 .SEQ_MODE=4'b1010;
    defparam \IR.ff8.q_0_fast_LC_2_14_7 .LUT_INIT=16'b1010111110100000;
    LogicCell40 \IR.ff8.q_0_fast_LC_2_14_7  (
            .in0(N__4387),
            .in1(_gnd_net_),
            .in2(N__8685),
            .in3(N__5291),
            .lcout(ir_out_fast_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVseq.counter.T_0_fast_2C_net ),
            .ce(),
            .sr(N__7304));
    defparam \IR.ff7.q_0_ner_LC_2_15_0 .C_ON=1'b0;
    defparam \IR.ff7.q_0_ner_LC_2_15_0 .SEQ_MODE=4'b1010;
    defparam \IR.ff7.q_0_ner_LC_2_15_0 .LUT_INIT=16'b1111111111110001;
    LogicCell40 \IR.ff7.q_0_ner_LC_2_15_0  (
            .in0(N__6525),
            .in1(N__6745),
            .in2(N__6836),
            .in3(N__6791),
            .lcout(ir_out_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVIR.ff7.q_0_nerC_net ),
            .ce(N__8687),
            .sr(N__7307));
    defparam \IR.ff6.q_0_ner_LC_2_15_1 .C_ON=1'b0;
    defparam \IR.ff6.q_0_ner_LC_2_15_1 .SEQ_MODE=4'b1010;
    defparam \IR.ff6.q_0_ner_LC_2_15_1 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \IR.ff6.q_0_ner_LC_2_15_1  (
            .in0(N__6692),
            .in1(N__6641),
            .in2(N__6605),
            .in3(N__6524),
            .lcout(ir_out_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVIR.ff7.q_0_nerC_net ),
            .ce(N__8687),
            .sr(N__7307));
    defparam \IR.ff8.q_0_ner_LC_2_15_2 .C_ON=1'b0;
    defparam \IR.ff8.q_0_ner_LC_2_15_2 .SEQ_MODE=4'b1010;
    defparam \IR.ff8.q_0_ner_LC_2_15_2 .LUT_INIT=16'b1111111111110001;
    LogicCell40 \IR.ff8.q_0_ner_LC_2_15_2  (
            .in0(N__6526),
            .in1(N__6900),
            .in2(N__6309),
            .in3(N__6334),
            .lcout(ir_out_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVIR.ff7.q_0_nerC_net ),
            .ce(N__8687),
            .sr(N__7307));
    defparam \seq.S0_0_i_N_3L3_LC_2_15_3 .C_ON=1'b0;
    defparam \seq.S0_0_i_N_3L3_LC_2_15_3 .SEQ_MODE=4'b0000;
    defparam \seq.S0_0_i_N_3L3_LC_2_15_3 .LUT_INIT=16'b0011001100000000;
    LogicCell40 \seq.S0_0_i_N_3L3_LC_2_15_3  (
            .in0(_gnd_net_),
            .in1(N__5281),
            .in2(_gnd_net_),
            .in3(N__3375),
            .lcout(\seq.S0_0_i_N_3LZ0Z3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.un1_ALU_en_0_1_LC_2_15_4 .C_ON=1'b0;
    defparam \seq.un1_ALU_en_0_1_LC_2_15_4 .SEQ_MODE=4'b0000;
    defparam \seq.un1_ALU_en_0_1_LC_2_15_4 .LUT_INIT=16'b0000101000001010;
    LogicCell40 \seq.un1_ALU_en_0_1_LC_2_15_4  (
            .in0(N__3376),
            .in1(_gnd_net_),
            .in2(N__5299),
            .in3(_gnd_net_),
            .lcout(\seq.un1_ALU_en_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \IR.ff4.q_ner_LC_2_15_6 .C_ON=1'b0;
    defparam \IR.ff4.q_ner_LC_2_15_6 .SEQ_MODE=4'b1010;
    defparam \IR.ff4.q_ner_LC_2_15_6 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \IR.ff4.q_ner_LC_2_15_6  (
            .in0(N__7740),
            .in1(N__7681),
            .in2(N__7593),
            .in3(N__7545),
            .lcout(ir_out_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVIR.ff7.q_0_nerC_net ),
            .ce(N__8687),
            .sr(N__7307));
    defparam \seq.counter.T_0_fast_RNIOL5V_2_LC_2_16_0 .C_ON=1'b0;
    defparam \seq.counter.T_0_fast_RNIOL5V_2_LC_2_16_0 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_0_fast_RNIOL5V_2_LC_2_16_0 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \seq.counter.T_0_fast_RNIOL5V_2_LC_2_16_0  (
            .in0(N__3356),
            .in1(N__4412),
            .in2(_gnd_net_),
            .in3(N__5547),
            .lcout(seq_un1_AR_OE_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.tbuf.g2_LC_2_16_1 .C_ON=1'b0;
    defparam \pc.tbuf.g2_LC_2_16_1 .SEQ_MODE=4'b0000;
    defparam \pc.tbuf.g2_LC_2_16_1 .LUT_INIT=16'b1101110101010101;
    LogicCell40 \pc.tbuf.g2_LC_2_16_1  (
            .in0(N__3875),
            .in1(N__3335),
            .in2(_gnd_net_),
            .in3(N__4587),
            .lcout(\pc.tbuf.gZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \AR.ff4.q_RNIT1RE_LC_2_16_3 .C_ON=1'b0;
    defparam \AR.ff4.q_RNIT1RE_LC_2_16_3 .SEQ_MODE=4'b0000;
    defparam \AR.ff4.q_RNIT1RE_LC_2_16_3 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \AR.ff4.q_RNIT1RE_LC_2_16_3  (
            .in0(N__3963),
            .in1(N__3926),
            .in2(_gnd_net_),
            .in3(N__5295),
            .lcout(),
            .ltout(g0_0_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.tbuf.g0_1_LC_2_16_4 .C_ON=1'b0;
    defparam \pc.tbuf.g0_1_LC_2_16_4 .SEQ_MODE=4'b0000;
    defparam \pc.tbuf.g0_1_LC_2_16_4 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \pc.tbuf.g0_1_LC_2_16_4  (
            .in0(N__3985),
            .in1(N__5827),
            .in2(N__3479),
            .in3(N__7400),
            .lcout(\pc.tbuf.g0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_RNIUILR_4_LC_2_16_6 .C_ON=1'b0;
    defparam \seq.counter.T_RNIUILR_4_LC_2_16_6 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_RNIUILR_4_LC_2_16_6 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \seq.counter.T_RNIUILR_4_LC_2_16_6  (
            .in0(N__5325),
            .in1(N__4411),
            .in2(_gnd_net_),
            .in3(N__5546),
            .lcout(\seq.counter.un7_ACC_LD_0 ),
            .ltout(\seq.counter.un7_ACC_LD_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_RNIK9TB2_4_LC_2_16_7 .C_ON=1'b0;
    defparam \seq.counter.T_RNIK9TB2_4_LC_2_16_7 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_RNIK9TB2_4_LC_2_16_7 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \seq.counter.T_RNIK9TB2_4_LC_2_16_7  (
            .in0(N__3467),
            .in1(N__5326),
            .in2(N__3461),
            .in3(N__5088),
            .lcout(seq_un1_ALU_en_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_0_RNILSL08_1_2_LC_4_8_1 .C_ON=1'b0;
    defparam \seq.counter.T_0_RNILSL08_1_2_LC_4_8_1 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_0_RNILSL08_1_2_LC_4_8_1 .LUT_INIT=16'b1100010000000000;
    LogicCell40 \seq.counter.T_0_RNILSL08_1_2_LC_4_8_1  (
            .in0(N__4667),
            .in1(N__4589),
            .in2(N__4943),
            .in3(N__4502),
            .lcout(IR_OE_2),
            .ltout(IR_OE_2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.tbuf.g0_8_LC_4_8_2 .C_ON=1'b0;
    defparam \pc.tbuf.g0_8_LC_4_8_2 .SEQ_MODE=4'b0000;
    defparam \pc.tbuf.g0_8_LC_4_8_2 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \pc.tbuf.g0_8_LC_4_8_2  (
            .in0(N__8435),
            .in1(N__8448),
            .in2(N__3458),
            .in3(N__8279),
            .lcout(bus_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_0_1_LC_4_9_0 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_0_1_LC_4_9_0 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_0_1_LC_4_9_0 .LUT_INIT=16'b1111111101111000;
    LogicCell40 \pc.program_counter_RNO_0_1_LC_4_9_0  (
            .in0(N__3670),
            .in1(N__8553),
            .in2(N__4838),
            .in3(N__3599),
            .lcout(\pc.program_counter_4_rn_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.un1_inc_LC_4_9_1 .C_ON=1'b0;
    defparam \pc.un1_inc_LC_4_9_1 .SEQ_MODE=4'b0000;
    defparam \pc.un1_inc_LC_4_9_1 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \pc.un1_inc_LC_4_9_1  (
            .in0(N__8552),
            .in1(N__4578),
            .in2(_gnd_net_),
            .in3(N__4213),
            .lcout(\pc.un1_inc_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_4_3_LC_4_9_4 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_4_3_LC_4_9_4 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_4_3_LC_4_9_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \pc.program_counter_RNO_4_3_LC_4_9_4  (
            .in0(_gnd_net_),
            .in1(N__3704),
            .in2(_gnd_net_),
            .in3(N__4832),
            .lcout(\pc.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_0_RNILSL08_2_LC_4_9_5 .C_ON=1'b0;
    defparam \seq.counter.T_0_RNILSL08_2_LC_4_9_5 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_0_RNILSL08_2_LC_4_9_5 .LUT_INIT=16'b1000110000000000;
    LogicCell40 \seq.counter.T_0_RNILSL08_2_LC_4_9_5  (
            .in0(N__3446),
            .in1(N__4577),
            .in2(N__4686),
            .in3(N__4492),
            .lcout(IR_OE_1),
            .ltout(IR_OE_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_1_1_LC_4_9_6 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_1_1_LC_4_9_6 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_1_1_LC_4_9_6 .LUT_INIT=16'b1111001100000000;
    LogicCell40 \pc.program_counter_RNO_1_1_LC_4_9_6  (
            .in0(_gnd_net_),
            .in1(N__8114),
            .in2(N__3602),
            .in3(N__3598),
            .lcout(\pc.program_counter_4_sn_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_RNIAFFM9_4_LC_4_9_7 .C_ON=1'b0;
    defparam \seq.counter.T_RNIAFFM9_4_LC_4_9_7 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_RNIAFFM9_4_LC_4_9_7 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \seq.counter.T_RNIAFFM9_4_LC_4_9_7  (
            .in0(N__5761),
            .in1(N__3731),
            .in2(N__5684),
            .in3(N__3824),
            .lcout(alu_out_m_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_2_0_LC_4_10_0 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_2_0_LC_4_10_0 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_2_0_LC_4_10_0 .LUT_INIT=16'b0000010001000100;
    LogicCell40 \pc.program_counter_RNO_2_0_LC_4_10_0  (
            .in0(N__4580),
            .in1(N__3578),
            .in2(N__4694),
            .in3(N__4267),
            .lcout(\pc.G_12_i_a3_2_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_6_0_LC_4_10_1 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_6_0_LC_4_10_1 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_6_0_LC_4_10_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \pc.program_counter_RNO_6_0_LC_4_10_1  (
            .in0(N__8549),
            .in1(N__8756),
            .in2(_gnd_net_),
            .in3(N__3514),
            .lcout(\pc.G_12_i_a3_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_RNO_0_0_LC_4_10_2 .C_ON=1'b0;
    defparam \seq.counter.T_RNO_0_0_LC_4_10_2 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_RNO_0_0_LC_4_10_2 .LUT_INIT=16'b0000000001010101;
    LogicCell40 \seq.counter.T_RNO_0_0_LC_4_10_2  (
            .in0(N__3515),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5188),
            .lcout(),
            .ltout(\seq.counter.T8_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_0_LC_4_10_3 .C_ON=1'b0;
    defparam \seq.counter.T_0_LC_4_10_3 .SEQ_MODE=4'b1011;
    defparam \seq.counter.T_0_LC_4_10_3 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \seq.counter.T_0_LC_4_10_3  (
            .in0(N__8551),
            .in1(N__4690),
            .in2(N__3572),
            .in3(N__5366),
            .lcout(seq_T_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVseq.counter.T_0C_net ),
            .ce(),
            .sr(N__7296));
    defparam \pc.program_counter_RNO_2_3_LC_4_10_4 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_2_3_LC_4_10_4 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_2_3_LC_4_10_4 .LUT_INIT=16'b0111111110000000;
    LogicCell40 \pc.program_counter_RNO_2_3_LC_4_10_4  (
            .in0(N__3662),
            .in1(N__8548),
            .in2(N__3569),
            .in3(N__4010),
            .lcout(\pc.N_188_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_1_LC_4_10_5 .C_ON=1'b0;
    defparam \seq.counter.T_1_LC_4_10_5 .SEQ_MODE=4'b1010;
    defparam \seq.counter.T_1_LC_4_10_5 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \seq.counter.T_1_LC_4_10_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3516),
            .lcout(inc),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVseq.counter.T_0C_net ),
            .ce(),
            .sr(N__7296));
    defparam \pc.program_counter_RNO_3_3_LC_4_10_7 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_3_3_LC_4_10_7 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_3_3_LC_4_10_7 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \pc.program_counter_RNO_3_3_LC_4_10_7  (
            .in0(N__8550),
            .in1(N__4579),
            .in2(_gnd_net_),
            .in3(N__4206),
            .lcout(\pc.un1_inc_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_1_2_LC_4_11_0 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_1_2_LC_4_11_0 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_1_2_LC_4_11_0 .LUT_INIT=16'b0100011100000011;
    LogicCell40 \pc.program_counter_RNO_1_2_LC_4_11_0  (
            .in0(N__5760),
            .in1(N__5679),
            .in2(N__3740),
            .in3(N__3820),
            .lcout(),
            .ltout(\pc.G_10_0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_2_LC_4_11_1 .C_ON=1'b0;
    defparam \pc.program_counter_2_LC_4_11_1 .SEQ_MODE=4'b1010;
    defparam \pc.program_counter_2_LC_4_11_1 .LUT_INIT=16'b1111111111101010;
    LogicCell40 \pc.program_counter_2_LC_4_11_1  (
            .in0(N__4088),
            .in1(N__3773),
            .in2(N__3752),
            .in3(N__3749),
            .lcout(\pc.program_counterZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4786),
            .ce(),
            .sr(N__7300));
    defparam \pc.program_counter_RNO_5_2_LC_4_11_2 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_5_2_LC_4_11_2 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_5_2_LC_4_11_2 .LUT_INIT=16'b0101101010101111;
    LogicCell40 \pc.program_counter_RNO_5_2_LC_4_11_2  (
            .in0(N__6162),
            .in1(_gnd_net_),
            .in2(N__8258),
            .in3(N__5990),
            .lcout(\pc.G_10_0_5_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.g0_3_LC_4_11_3 .C_ON=1'b0;
    defparam \ALU_main.g0_3_LC_4_11_3 .SEQ_MODE=4'b0000;
    defparam \ALU_main.g0_3_LC_4_11_3 .LUT_INIT=16'b1000100001100110;
    LogicCell40 \ALU_main.g0_3_LC_4_11_3  (
            .in0(N__5991),
            .in1(N__8257),
            .in2(_gnd_net_),
            .in3(N__6163),
            .lcout(ALU_main_N_43_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.un1_A_axb_2_l_ofx_LC_4_11_5 .C_ON=1'b0;
    defparam \ALU_main.un1_A_axb_2_l_ofx_LC_4_11_5 .SEQ_MODE=4'b0000;
    defparam \ALU_main.un1_A_axb_2_l_ofx_LC_4_11_5 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU_main.un1_A_axb_2_l_ofx_LC_4_11_5  (
            .in0(N__5992),
            .in1(N__8253),
            .in2(_gnd_net_),
            .in3(N__6161),
            .lcout(\ALU_main.un1_A_axb_2_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_4_2_LC_4_11_7 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_4_2_LC_4_11_7 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_4_2_LC_4_11_7 .LUT_INIT=16'b0110011011001100;
    LogicCell40 \pc.program_counter_RNO_4_2_LC_4_11_7  (
            .in0(N__4833),
            .in1(N__3700),
            .in2(_gnd_net_),
            .in3(N__3666),
            .lcout(\pc.N_10_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.un1_A_cry_0_c_THRU_CRY_0_LC_4_12_0 .C_ON=1'b1;
    defparam \ALU_main.un1_A_cry_0_c_THRU_CRY_0_LC_4_12_0 .SEQ_MODE=4'b0000;
    defparam \ALU_main.un1_A_cry_0_c_THRU_CRY_0_LC_4_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \ALU_main.un1_A_cry_0_c_THRU_CRY_0_LC_4_12_0  (
            .in0(_gnd_net_),
            .in1(N__3622),
            .in2(N__3626),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_12_0_),
            .carryout(\ALU_main.un1_A_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.un1_A_cry_0_s_LC_4_12_1 .C_ON=1'b1;
    defparam \ALU_main.un1_A_cry_0_s_LC_4_12_1 .SEQ_MODE=4'b0000;
    defparam \ALU_main.un1_A_cry_0_s_LC_4_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU_main.un1_A_cry_0_s_LC_4_12_1  (
            .in0(_gnd_net_),
            .in1(N__6060),
            .in2(N__4928),
            .in3(N__3608),
            .lcout(un1_A_cry_0_s),
            .ltout(),
            .carryin(\ALU_main.un1_A_cry_0_c_THRU_CO ),
            .carryout(\ALU_main.un1_A_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.un1_A_cry_0_c_RNIPCLO2_LC_4_12_2 .C_ON=1'b1;
    defparam \ALU_main.un1_A_cry_0_c_RNIPCLO2_LC_4_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU_main.un1_A_cry_0_c_RNIPCLO2_LC_4_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU_main.un1_A_cry_0_c_RNIPCLO2_LC_4_12_2  (
            .in0(_gnd_net_),
            .in1(N__6028),
            .in2(N__5060),
            .in3(N__3605),
            .lcout(un1_A_cry_0_c_RNIPCLO2),
            .ltout(),
            .carryin(\ALU_main.un1_A_cry_0 ),
            .carryout(\ALU_main.un1_A_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.un1_A_cry_1_c_RNITKPO2_LC_4_12_3 .C_ON=1'b1;
    defparam \ALU_main.un1_A_cry_1_c_RNITKPO2_LC_4_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU_main.un1_A_cry_1_c_RNITKPO2_LC_4_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU_main.un1_A_cry_1_c_RNITKPO2_LC_4_12_3  (
            .in0(_gnd_net_),
            .in1(N__5989),
            .in2(N__3833),
            .in3(N__3809),
            .lcout(un1_A_cry_1_c_RNITKPO2),
            .ltout(),
            .carryin(\ALU_main.un1_A_cry_1 ),
            .carryout(\ALU_main.un1_A_cry_2 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.un1_A_cry_2_c_RNI1TTO2_LC_4_12_4 .C_ON=1'b1;
    defparam \ALU_main.un1_A_cry_2_c_RNI1TTO2_LC_4_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU_main.un1_A_cry_2_c_RNI1TTO2_LC_4_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU_main.un1_A_cry_2_c_RNI1TTO2_LC_4_12_4  (
            .in0(_gnd_net_),
            .in1(N__4919),
            .in2(N__5828),
            .in3(N__3806),
            .lcout(un1_A_cry_2_c_RNI1TTO2),
            .ltout(),
            .carryin(\ALU_main.un1_A_cry_2 ),
            .carryout(\ALU_main.un1_A_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.un1_A_cry_3_c_RNI552P2_LC_4_12_5 .C_ON=1'b1;
    defparam \ALU_main.un1_A_cry_3_c_RNI552P2_LC_4_12_5 .SEQ_MODE=4'b0000;
    defparam \ALU_main.un1_A_cry_3_c_RNI552P2_LC_4_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU_main.un1_A_cry_3_c_RNI552P2_LC_4_12_5  (
            .in0(_gnd_net_),
            .in1(N__5051),
            .in2(N__7908),
            .in3(N__3803),
            .lcout(\ALU_main.un1_A_cry_3_c_RNI552PZ0Z2 ),
            .ltout(),
            .carryin(\ALU_main.un1_A_cry_3 ),
            .carryout(\ALU_main.un1_A_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.un1_A_cry_4_c_RNI9D6P2_LC_4_12_6 .C_ON=1'b1;
    defparam \ALU_main.un1_A_cry_4_c_RNI9D6P2_LC_4_12_6 .SEQ_MODE=4'b0000;
    defparam \ALU_main.un1_A_cry_4_c_RNI9D6P2_LC_4_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU_main.un1_A_cry_4_c_RNI9D6P2_LC_4_12_6  (
            .in0(_gnd_net_),
            .in1(N__5228),
            .in2(N__5855),
            .in3(N__3800),
            .lcout(\ALU_main.un1_A_cry_4_c_RNI9D6PZ0Z2 ),
            .ltout(),
            .carryin(\ALU_main.un1_A_cry_4 ),
            .carryout(\ALU_main.un1_A_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.un1_A_cry_5_c_RNIDLAP2_LC_4_12_7 .C_ON=1'b1;
    defparam \ALU_main.un1_A_cry_5_c_RNIDLAP2_LC_4_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU_main.un1_A_cry_5_c_RNIDLAP2_LC_4_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \ALU_main.un1_A_cry_5_c_RNIDLAP2_LC_4_12_7  (
            .in0(_gnd_net_),
            .in1(N__5885),
            .in2(N__5912),
            .in3(N__3797),
            .lcout(\ALU_main.un1_A_cry_5_c_RNIDLAPZ0Z2 ),
            .ltout(),
            .carryin(\ALU_main.un1_A_cry_5 ),
            .carryout(\ALU_main.un1_A_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.un1_A_cry_6_c_RNIP89E2_LC_4_13_0 .C_ON=1'b0;
    defparam \ALU_main.un1_A_cry_6_c_RNIP89E2_LC_4_13_0 .SEQ_MODE=4'b0000;
    defparam \ALU_main.un1_A_cry_6_c_RNIP89E2_LC_4_13_0 .LUT_INIT=16'b1001011001101001;
    LogicCell40 \ALU_main.un1_A_cry_6_c_RNIP89E2_LC_4_13_0  (
            .in0(N__6167),
            .in1(N__5866),
            .in2(N__6268),
            .in3(N__3794),
            .lcout(\ALU_main.un1_A_cry_6_c_RNIP89EZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \mem.data_2_7_0__g0_1_LC_4_13_1 .C_ON=1'b0;
    defparam \mem.data_2_7_0__g0_1_LC_4_13_1 .SEQ_MODE=4'b0000;
    defparam \mem.data_2_7_0__g0_1_LC_4_13_1 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \mem.data_2_7_0__g0_1_LC_4_13_1  (
            .in0(N__4118),
            .in1(N__5748),
            .in2(N__4079),
            .in3(N__5675),
            .lcout(alu_out_m_1_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.un1_A_cry_5_c_RNI209N9_LC_4_13_2 .C_ON=1'b0;
    defparam \ALU_main.un1_A_cry_5_c_RNI209N9_LC_4_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU_main.un1_A_cry_5_c_RNI209N9_LC_4_13_2 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \ALU_main.un1_A_cry_5_c_RNI209N9_LC_4_13_2  (
            .in0(N__5747),
            .in1(N__3779),
            .in2(N__5924),
            .in3(N__5674),
            .lcout(alu_out_m_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.g0_LC_4_13_3 .C_ON=1'b0;
    defparam \ALU_main.g0_LC_4_13_3 .SEQ_MODE=4'b0000;
    defparam \ALU_main.g0_LC_4_13_3 .LUT_INIT=16'b1000100001100110;
    LogicCell40 \ALU_main.g0_LC_4_13_3  (
            .in0(N__5820),
            .in1(N__7833),
            .in2(_gnd_net_),
            .in3(N__6166),
            .lcout(),
            .ltout(ALU_main_N_44_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \mem.data_2_7_0__g0_0_LC_4_13_4 .C_ON=1'b0;
    defparam \mem.data_2_7_0__g0_0_LC_4_13_4 .SEQ_MODE=4'b0000;
    defparam \mem.data_2_7_0__g0_0_LC_4_13_4 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \mem.data_2_7_0__g0_0_LC_4_13_4  (
            .in0(N__5746),
            .in1(N__5673),
            .in2(N__4121),
            .in3(N__4117),
            .lcout(alu_out_m_0_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_0_2_LC_4_13_6 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_0_2_LC_4_13_6 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_0_2_LC_4_13_6 .LUT_INIT=16'b1101100010001000;
    LogicCell40 \pc.program_counter_RNO_0_2_LC_4_13_6  (
            .in0(N__8621),
            .in1(N__4109),
            .in2(N__8434),
            .in3(N__4100),
            .lcout(\pc.G_10_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.g0_0_LC_4_13_7 .C_ON=1'b0;
    defparam \ALU_main.g0_0_LC_4_13_7 .SEQ_MODE=4'b0000;
    defparam \ALU_main.g0_0_LC_4_13_7 .LUT_INIT=16'b1000100001100110;
    LogicCell40 \ALU_main.g0_0_LC_4_13_7  (
            .in0(N__5821),
            .in1(N__7834),
            .in2(_gnd_net_),
            .in3(N__6168),
            .lcout(ALU_main_N_44_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.tbuf.g0_0_1_LC_4_14_1 .C_ON=1'b0;
    defparam \pc.tbuf.g0_0_1_LC_4_14_1 .SEQ_MODE=4'b0000;
    defparam \pc.tbuf.g0_0_1_LC_4_14_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \pc.tbuf.g0_0_1_LC_4_14_1  (
            .in0(_gnd_net_),
            .in1(N__5823),
            .in2(_gnd_net_),
            .in3(N__7412),
            .lcout(\pc.tbuf.g0_0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_1_3_LC_4_14_2 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_1_3_LC_4_14_2 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_1_3_LC_4_14_2 .LUT_INIT=16'b1000100010000000;
    LogicCell40 \pc.program_counter_RNO_1_3_LC_4_14_2  (
            .in0(N__4070),
            .in1(N__4061),
            .in2(N__4049),
            .in3(N__6527),
            .lcout(),
            .ltout(\pc.g0_sn_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_3_LC_4_14_3 .C_ON=1'b0;
    defparam \pc.program_counter_3_LC_4_14_3 .SEQ_MODE=4'b1010;
    defparam \pc.program_counter_3_LC_4_14_3 .LUT_INIT=16'b1111101011001010;
    LogicCell40 \pc.program_counter_3_LC_4_14_3  (
            .in0(N__4031),
            .in1(N__3839),
            .in2(N__4019),
            .in3(N__4016),
            .lcout(\pc.program_counterZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4796),
            .ce(),
            .sr(N__7310));
    defparam \AR.ff4.q_RNILN0E1_LC_4_14_4 .C_ON=1'b0;
    defparam \AR.ff4.q_RNILN0E1_LC_4_14_4 .SEQ_MODE=4'b0000;
    defparam \AR.ff4.q_RNILN0E1_LC_4_14_4 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \AR.ff4.q_RNILN0E1_LC_4_14_4  (
            .in0(N__3989),
            .in1(N__3971),
            .in2(N__3925),
            .in3(N__5312),
            .lcout(),
            .ltout(AR_out_m_3_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.tbuf.g0_0_LC_4_14_5 .C_ON=1'b0;
    defparam \pc.tbuf.g0_0_LC_4_14_5 .SEQ_MODE=4'b0000;
    defparam \pc.tbuf.g0_0_LC_4_14_5 .LUT_INIT=16'b1111001111111011;
    LogicCell40 \pc.tbuf.g0_0_LC_4_14_5  (
            .in0(N__3889),
            .in1(N__3848),
            .in2(N__3842),
            .in3(N__4493),
            .lcout(\pc.g0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \IR.ff6.q_0_ner_RNIVL0RI_LC_4_15_1 .C_ON=1'b0;
    defparam \IR.ff6.q_0_ner_RNIVL0RI_LC_4_15_1 .SEQ_MODE=4'b0000;
    defparam \IR.ff6.q_0_ner_RNIVL0RI_LC_4_15_1 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \IR.ff6.q_0_ner_RNIVL0RI_LC_4_15_1  (
            .in0(N__8673),
            .in1(N__6079),
            .in2(_gnd_net_),
            .in3(N__4418),
            .lcout(N_2_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \IR.ff8.q_0_ner_RNIND22I_LC_4_15_2 .C_ON=1'b0;
    defparam \IR.ff8.q_0_ner_RNIND22I_LC_4_15_2 .SEQ_MODE=4'b0000;
    defparam \IR.ff8.q_0_ner_RNIND22I_LC_4_15_2 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \IR.ff8.q_0_ner_RNIND22I_LC_4_15_2  (
            .in0(N__8677),
            .in1(N__4388),
            .in2(_gnd_net_),
            .in3(N__5309),
            .lcout(),
            .ltout(N_1_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.q_ret_1_LC_4_15_3 .C_ON=1'b0;
    defparam \seq.q_ret_1_LC_4_15_3 .SEQ_MODE=4'b1010;
    defparam \seq.q_ret_1_LC_4_15_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \seq.q_ret_1_LC_4_15_3  (
            .in0(N__5510),
            .in1(N__4358),
            .in2(N__4340),
            .in3(N__4322),
            .lcout(seq_un1_HLT_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVseq.q_ret_1C_net ),
            .ce(),
            .sr(N__7314));
    defparam \seq.counter.T_RNI1G50J_1_LC_4_15_4 .C_ON=1'b0;
    defparam \seq.counter.T_RNI1G50J_1_LC_4_15_4 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_RNI1G50J_1_LC_4_15_4 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \seq.counter.T_RNI1G50J_1_LC_4_15_4  (
            .in0(_gnd_net_),
            .in1(N__8674),
            .in2(_gnd_net_),
            .in3(N__4308),
            .lcout(\seq.un1_HLT_1_reti ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.q_ret_LC_4_16_5 .C_ON=1'b0;
    defparam \seq.q_ret_LC_4_16_5 .SEQ_MODE=4'b1010;
    defparam \seq.q_ret_LC_4_16_5 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \seq.q_ret_LC_4_16_5  (
            .in0(_gnd_net_),
            .in1(N__8675),
            .in2(_gnd_net_),
            .in3(N__4309),
            .lcout(\seq.un1_HLT_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVseq.q_retC_net ),
            .ce(),
            .sr(N__7319));
    defparam \pc.tbuf.g0_6_LC_5_9_0 .C_ON=1'b0;
    defparam \pc.tbuf.g0_6_LC_5_9_0 .SEQ_MODE=4'b0000;
    defparam \pc.tbuf.g0_6_LC_5_9_0 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \pc.tbuf.g0_6_LC_5_9_0  (
            .in0(N__8166),
            .in1(N__8210),
            .in2(N__8129),
            .in3(N__8060),
            .lcout(),
            .ltout(bus_1_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \AR.ff2.q_LC_5_9_1 .C_ON=1'b0;
    defparam \AR.ff2.q_LC_5_9_1 .SEQ_MODE=4'b1010;
    defparam \AR.ff2.q_LC_5_9_1 .LUT_INIT=16'b1110001010101010;
    LogicCell40 \AR.ff2.q_LC_5_9_1  (
            .in0(N__4135),
            .in1(N__4692),
            .in2(N__4277),
            .in3(N__4274),
            .lcout(AR_out_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVAR.ff2.qC_net ),
            .ce(),
            .sr(N__7293));
    defparam \pc.tbuf.out_1_1_iv_0_LC_5_9_2 .C_ON=1'b0;
    defparam \pc.tbuf.out_1_1_iv_0_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \pc.tbuf.out_1_1_iv_0_LC_5_9_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \pc.tbuf.out_1_1_iv_0_LC_5_9_2  (
            .in0(N__6024),
            .in1(N__4214),
            .in2(N__4136),
            .in3(N__7476),
            .lcout(\pc.tbuf.out_1_1_ivZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_3_LC_5_9_3 .C_ON=1'b0;
    defparam \seq.counter.T_3_LC_5_9_3 .SEQ_MODE=4'b1010;
    defparam \seq.counter.T_3_LC_5_9_3 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \seq.counter.T_3_LC_5_9_3  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__4693),
            .lcout(\seq.counter.TZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVAR.ff2.qC_net ),
            .ce(),
            .sr(N__7293));
    defparam \seq.counter.T_RNIPO8O2_3_LC_5_9_5 .C_ON=1'b0;
    defparam \seq.counter.T_RNIPO8O2_3_LC_5_9_5 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_RNIPO8O2_3_LC_5_9_5 .LUT_INIT=16'b0001001101011111;
    LogicCell40 \seq.counter.T_RNIPO8O2_3_LC_5_9_5  (
            .in0(N__4982),
            .in1(N__5096),
            .in2(N__5202),
            .in3(N__5364),
            .lcout(),
            .ltout(\seq.counter.ACC_LD_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_RNIIRQM5_4_LC_5_9_6 .C_ON=1'b0;
    defparam \seq.counter.T_RNIIRQM5_4_LC_5_9_6 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_RNIIRQM5_4_LC_5_9_6 .LUT_INIT=16'b1000111111111111;
    LogicCell40 \seq.counter.T_RNIIRQM5_4_LC_5_9_6  (
            .in0(N__5365),
            .in1(N__4904),
            .in2(N__4874),
            .in3(N__6193),
            .lcout(seq_ACC_LD_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \mem.data_2_7_0__g0_i_LC_5_10_3 .C_ON=1'b0;
    defparam \mem.data_2_7_0__g0_i_LC_5_10_3 .SEQ_MODE=4'b0000;
    defparam \mem.data_2_7_0__g0_i_LC_5_10_3 .LUT_INIT=16'b0111101111001111;
    LogicCell40 \mem.data_2_7_0__g0_i_LC_5_10_3  (
            .in0(N__7167),
            .in1(N__7108),
            .in2(N__7053),
            .in3(N__6968),
            .lcout(),
            .ltout(mem_data_2_7_0__N_11_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.tbuf.g0_7_LC_5_10_4 .C_ON=1'b0;
    defparam \pc.tbuf.g0_7_LC_5_10_4 .SEQ_MODE=4'b0000;
    defparam \pc.tbuf.g0_7_LC_5_10_4 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \pc.tbuf.g0_7_LC_5_10_4  (
            .in0(N__4871),
            .in1(N__4862),
            .in2(N__4856),
            .in3(N__6537),
            .lcout(\pc.g0_1_0 ),
            .ltout(\pc.g0_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_1_LC_5_10_5 .C_ON=1'b0;
    defparam \pc.program_counter_1_LC_5_10_5 .SEQ_MODE=4'b1010;
    defparam \pc.program_counter_1_LC_5_10_5 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \pc.program_counter_1_LC_5_10_5  (
            .in0(N__4853),
            .in1(N__4847),
            .in2(N__4841),
            .in3(N__8045),
            .lcout(\pc.program_counterZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__4787),
            .ce(),
            .sr(N__7301));
    defparam \seq.counter.T_0_RNILSL08_0_2_LC_5_11_0 .C_ON=1'b0;
    defparam \seq.counter.T_0_RNILSL08_0_2_LC_5_11_0 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_0_RNILSL08_0_2_LC_5_11_0 .LUT_INIT=16'b1100010000000000;
    LogicCell40 \seq.counter.T_0_RNILSL08_0_2_LC_5_11_0  (
            .in0(N__4691),
            .in1(N__4588),
            .in2(N__4430),
            .in3(N__4501),
            .lcout(IR_OE_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.g2_LC_5_11_1 .C_ON=1'b0;
    defparam \seq.g2_LC_5_11_1 .SEQ_MODE=4'b0000;
    defparam \seq.g2_LC_5_11_1 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \seq.g2_LC_5_11_1  (
            .in0(N__4980),
            .in1(N__5155),
            .in2(_gnd_net_),
            .in3(N__5014),
            .lcout(\seq.gZ0Z2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.g0_2_LC_5_11_2 .C_ON=1'b0;
    defparam \ALU_main.g0_2_LC_5_11_2 .SEQ_MODE=4'b0000;
    defparam \ALU_main.g0_2_LC_5_11_2 .LUT_INIT=16'b1001100101000100;
    LogicCell40 \ALU_main.g0_2_LC_5_11_2  (
            .in0(N__6157),
            .in1(N__6014),
            .in2(_gnd_net_),
            .in3(N__6854),
            .lcout(),
            .ltout(ALU_main_N_42_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_RNI439M9_4_LC_5_11_3 .C_ON=1'b0;
    defparam \seq.counter.T_RNI439M9_4_LC_5_11_3 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_RNI439M9_4_LC_5_11_3 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \seq.counter.T_RNI439M9_4_LC_5_11_3  (
            .in0(N__5762),
            .in1(N__5682),
            .in2(N__5045),
            .in3(N__5042),
            .lcout(alu_out_m_0_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.g0_1_LC_5_11_4 .C_ON=1'b0;
    defparam \ALU_main.g0_1_LC_5_11_4 .SEQ_MODE=4'b0000;
    defparam \ALU_main.g0_1_LC_5_11_4 .LUT_INIT=16'b1001100101000100;
    LogicCell40 \ALU_main.g0_1_LC_5_11_4  (
            .in0(N__6158),
            .in1(N__6050),
            .in2(_gnd_net_),
            .in3(N__6244),
            .lcout(),
            .ltout(ALU_main_N_41_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_RNIP3LPB_4_LC_5_11_5 .C_ON=1'b0;
    defparam \seq.counter.T_RNIP3LPB_4_LC_5_11_5 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_RNIP3LPB_4_LC_5_11_5 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \seq.counter.T_RNIP3LPB_4_LC_5_11_5  (
            .in0(N__5763),
            .in1(N__5683),
            .in2(N__5036),
            .in3(N__5029),
            .lcout(alu_out_m_0_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.g2_1_LC_5_11_6 .C_ON=1'b0;
    defparam \seq.g2_1_LC_5_11_6 .SEQ_MODE=4'b0000;
    defparam \seq.g2_1_LC_5_11_6 .LUT_INIT=16'b0000000000010001;
    LogicCell40 \seq.g2_1_LC_5_11_6  (
            .in0(N__5015),
            .in1(N__4981),
            .in2(_gnd_net_),
            .in3(N__5156),
            .lcout(\seq.g2Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.un1_A_axb_0_l_ofx_LC_5_11_7 .C_ON=1'b0;
    defparam \ALU_main.un1_A_axb_0_l_ofx_LC_5_11_7 .SEQ_MODE=4'b0000;
    defparam \ALU_main.un1_A_axb_0_l_ofx_LC_5_11_7 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \ALU_main.un1_A_axb_0_l_ofx_LC_5_11_7  (
            .in0(N__6243),
            .in1(N__6051),
            .in2(_gnd_net_),
            .in3(N__6156),
            .lcout(\ALU_main.un1_A_axb_0_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \acc.ff6.q_RNI207H1_LC_5_12_0 .C_ON=1'b0;
    defparam \acc.ff6.q_RNI207H1_LC_5_12_0 .SEQ_MODE=4'b0000;
    defparam \acc.ff6.q_RNI207H1_LC_5_12_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \acc.ff6.q_RNI207H1_LC_5_12_0  (
            .in0(N__5853),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7454),
            .lcout(acc_out_m_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.un1_A_axb_3_l_ofx_LC_5_12_2 .C_ON=1'b0;
    defparam \ALU_main.un1_A_axb_3_l_ofx_LC_5_12_2 .SEQ_MODE=4'b0000;
    defparam \ALU_main.un1_A_axb_3_l_ofx_LC_5_12_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU_main.un1_A_axb_3_l_ofx_LC_5_12_2  (
            .in0(N__5822),
            .in1(N__7835),
            .in2(_gnd_net_),
            .in3(N__6164),
            .lcout(\ALU_main.un1_A_axb_3_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.ALU_Out_0_5_LC_5_12_3 .C_ON=1'b0;
    defparam \ALU_main.ALU_Out_0_5_LC_5_12_3 .SEQ_MODE=4'b0000;
    defparam \ALU_main.ALU_Out_0_5_LC_5_12_3 .LUT_INIT=16'b1001100101000100;
    LogicCell40 \ALU_main.ALU_Out_0_5_LC_5_12_3  (
            .in0(N__6165),
            .in1(N__5852),
            .in2(_gnd_net_),
            .in3(N__6359),
            .lcout(),
            .ltout(\ALU_main.N_46_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.un1_A_cry_4_c_RNISJ2N9_LC_5_12_4 .C_ON=1'b0;
    defparam \ALU_main.un1_A_cry_4_c_RNISJ2N9_LC_5_12_4 .SEQ_MODE=4'b0000;
    defparam \ALU_main.un1_A_cry_4_c_RNISJ2N9_LC_5_12_4 .LUT_INIT=16'b0100010011110000;
    LogicCell40 \ALU_main.un1_A_cry_4_c_RNISJ2N9_LC_5_12_4  (
            .in0(N__5768),
            .in1(N__4913),
            .in2(N__4907),
            .in3(N__5680),
            .lcout(alu_out_m_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.g0_i_a3_0_2_LC_5_12_5 .C_ON=1'b0;
    defparam \seq.g0_i_a3_0_2_LC_5_12_5 .SEQ_MODE=4'b0000;
    defparam \seq.g0_i_a3_0_2_LC_5_12_5 .LUT_INIT=16'b0010001000000000;
    LogicCell40 \seq.g0_i_a3_0_2_LC_5_12_5  (
            .in0(N__5504),
            .in1(N__5456),
            .in2(_gnd_net_),
            .in3(N__5406),
            .lcout(),
            .ltout(\seq.g0_i_a3_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_RNI51KH1_4_LC_5_12_6 .C_ON=1'b0;
    defparam \seq.counter.T_RNI51KH1_4_LC_5_12_6 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_RNI51KH1_4_LC_5_12_6 .LUT_INIT=16'b1101110111011111;
    LogicCell40 \seq.counter.T_RNI51KH1_4_LC_5_12_6  (
            .in0(N__5363),
            .in1(N__5310),
            .in2(N__5246),
            .in3(N__5243),
            .lcout(seq_S0_0),
            .ltout(seq_S0_0_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.un1_A_axb_5_l_ofx_LC_5_12_7 .C_ON=1'b0;
    defparam \ALU_main.un1_A_axb_5_l_ofx_LC_5_12_7 .SEQ_MODE=4'b0000;
    defparam \ALU_main.un1_A_axb_5_l_ofx_LC_5_12_7 .LUT_INIT=16'b1111000000001111;
    LogicCell40 \ALU_main.un1_A_axb_5_l_ofx_LC_5_12_7  (
            .in0(_gnd_net_),
            .in1(N__5854),
            .in2(N__5231),
            .in3(N__6358),
            .lcout(\ALU_main.un1_A_axb_5_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \seq.counter.T_RNIR83I4_3_LC_5_13_0 .C_ON=1'b0;
    defparam \seq.counter.T_RNIR83I4_3_LC_5_13_0 .SEQ_MODE=4'b0000;
    defparam \seq.counter.T_RNIR83I4_3_LC_5_13_0 .LUT_INIT=16'b1010101010001010;
    LogicCell40 \seq.counter.T_RNIR83I4_3_LC_5_13_0  (
            .in0(N__5203),
            .in1(N__5154),
            .in2(N__5108),
            .in3(N__5092),
            .lcout(seq_B_LD_0_i),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.un1_A_axb_1_l_ofx_LC_5_13_2 .C_ON=1'b0;
    defparam \ALU_main.un1_A_axb_1_l_ofx_LC_5_13_2 .SEQ_MODE=4'b0000;
    defparam \ALU_main.un1_A_axb_1_l_ofx_LC_5_13_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU_main.un1_A_axb_1_l_ofx_LC_5_13_2  (
            .in0(N__6029),
            .in1(N__6847),
            .in2(_gnd_net_),
            .in3(N__6159),
            .lcout(\ALU_main.un1_A_axb_1_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b_reg.ff5.q_LC_5_13_4 .C_ON=1'b0;
    defparam \b_reg.ff5.q_LC_5_13_4 .SEQ_MODE=4'b1010;
    defparam \b_reg.ff5.q_LC_5_13_4 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \b_reg.ff5.q_LC_5_13_4  (
            .in0(N__7951),
            .in1(N__7994),
            .in2(N__7914),
            .in3(N__7456),
            .lcout(b_reg_out_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVb_reg.ff5.qC_net ),
            .ce(N__7781),
            .sr(N__7311));
    defparam \ALU_main.un1_A_axb_4_l_ofx_LC_5_13_5 .C_ON=1'b0;
    defparam \ALU_main.un1_A_axb_4_l_ofx_LC_5_13_5 .SEQ_MODE=4'b0000;
    defparam \ALU_main.un1_A_axb_4_l_ofx_LC_5_13_5 .LUT_INIT=16'b1010101001010101;
    LogicCell40 \ALU_main.un1_A_axb_4_l_ofx_LC_5_13_5  (
            .in0(N__6160),
            .in1(N__7903),
            .in2(_gnd_net_),
            .in3(N__6205),
            .lcout(\ALU_main.un1_A_axb_4_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \acc.ff7.q_RNI328H1_LC_5_13_6 .C_ON=1'b0;
    defparam \acc.ff7.q_RNI328H1_LC_5_13_6 .SEQ_MODE=4'b0000;
    defparam \acc.ff7.q_RNI328H1_LC_5_13_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \acc.ff7.q_RNI328H1_LC_5_13_6  (
            .in0(_gnd_net_),
            .in1(N__5908),
            .in2(_gnd_net_),
            .in3(N__7455),
            .lcout(acc_out_m_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \acc.ff7.q_LC_5_14_0 .C_ON=1'b0;
    defparam \acc.ff7.q_LC_5_14_0 .SEQ_MODE=4'b1010;
    defparam \acc.ff7.q_LC_5_14_0 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \acc.ff7.q_LC_5_14_0  (
            .in0(N__6821),
            .in1(N__6778),
            .in2(N__6735),
            .in3(N__6535),
            .lcout(acc_out_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVacc.ff7.qC_net ),
            .ce(N__5948),
            .sr(N__7315));
    defparam \ALU_main.ALU_Out_0_6_LC_5_14_1 .C_ON=1'b0;
    defparam \ALU_main.ALU_Out_0_6_LC_5_14_1 .SEQ_MODE=4'b0000;
    defparam \ALU_main.ALU_Out_0_6_LC_5_14_1 .LUT_INIT=16'b1001100101000100;
    LogicCell40 \ALU_main.ALU_Out_0_6_LC_5_14_1  (
            .in0(N__6191),
            .in1(N__5906),
            .in2(_gnd_net_),
            .in3(N__6704),
            .lcout(\ALU_main.N_47 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.un1_A_axb_6_l_ofx_LC_5_14_2 .C_ON=1'b0;
    defparam \ALU_main.un1_A_axb_6_l_ofx_LC_5_14_2 .SEQ_MODE=4'b0000;
    defparam \ALU_main.un1_A_axb_6_l_ofx_LC_5_14_2 .LUT_INIT=16'b1100110000110011;
    LogicCell40 \ALU_main.un1_A_axb_6_l_ofx_LC_5_14_2  (
            .in0(N__5907),
            .in1(N__6703),
            .in2(_gnd_net_),
            .in3(N__6190),
            .lcout(\ALU_main.un1_A_axb_6_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \acc.ff8.q_LC_5_14_3 .C_ON=1'b0;
    defparam \acc.ff8.q_LC_5_14_3 .SEQ_MODE=4'b1010;
    defparam \acc.ff8.q_LC_5_14_3 .LUT_INIT=16'b1111111111001101;
    LogicCell40 \acc.ff8.q_LC_5_14_3  (
            .in0(N__6536),
            .in1(N__6350),
            .in2(N__6891),
            .in3(N__6310),
            .lcout(acc_out_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVacc.ff7.qC_net ),
            .ce(N__5948),
            .sr(N__7315));
    defparam \acc.ff6.q_LC_5_14_4 .C_ON=1'b0;
    defparam \acc.ff6.q_LC_5_14_4 .SEQ_MODE=4'b1010;
    defparam \acc.ff6.q_LC_5_14_4 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \acc.ff6.q_LC_5_14_4  (
            .in0(N__6636),
            .in1(N__6683),
            .in2(N__6599),
            .in3(N__6534),
            .lcout(acc_out_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVacc.ff7.qC_net ),
            .ce(N__5948),
            .sr(N__7315));
    defparam \acc.ff4.q_LC_5_14_6 .C_ON=1'b0;
    defparam \acc.ff4.q_LC_5_14_6 .SEQ_MODE=4'b1010;
    defparam \acc.ff4.q_LC_5_14_6 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \acc.ff4.q_LC_5_14_6  (
            .in0(N__7741),
            .in1(N__7680),
            .in2(N__7619),
            .in3(N__7524),
            .lcout(acc_out_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVacc.ff7.qC_net ),
            .ce(N__5948),
            .sr(N__7315));
    defparam \ALU_main.un1_A_cry_3_c_RNIM7SM9_LC_5_15_0 .C_ON=1'b0;
    defparam \ALU_main.un1_A_cry_3_c_RNIM7SM9_LC_5_15_0 .SEQ_MODE=4'b0000;
    defparam \ALU_main.un1_A_cry_3_c_RNIM7SM9_LC_5_15_0 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \ALU_main.un1_A_cry_3_c_RNIM7SM9_LC_5_15_0  (
            .in0(N__5777),
            .in1(N__5767),
            .in2(N__6095),
            .in3(N__5681),
            .lcout(alu_out_m_4),
            .ltout(alu_out_m_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buf1.out_1_2_iv_LC_5_15_1 .C_ON=1'b0;
    defparam \buf1.out_1_2_iv_LC_5_15_1 .SEQ_MODE=4'b0000;
    defparam \buf1.out_1_2_iv_LC_5_15_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \buf1.out_1_2_iv_LC_5_15_1  (
            .in0(N__7910),
            .in1(N__7959),
            .in2(N__5597),
            .in3(N__7457),
            .lcout(bus_4),
            .ltout(bus_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \IR.ff5.q_0_ner_RNINVSHI_LC_5_15_2 .C_ON=1'b0;
    defparam \IR.ff5.q_0_ner_RNINVSHI_LC_5_15_2 .SEQ_MODE=4'b0000;
    defparam \IR.ff5.q_0_ner_RNINVSHI_LC_5_15_2 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \IR.ff5.q_0_ner_RNINVSHI_LC_5_15_2  (
            .in0(_gnd_net_),
            .in1(N__8676),
            .in2(N__5567),
            .in3(N__5563),
            .lcout(N_4_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \ALU_main.ALU_Out_0_4_LC_5_15_5 .C_ON=1'b0;
    defparam \ALU_main.ALU_Out_0_4_LC_5_15_5 .SEQ_MODE=4'b0000;
    defparam \ALU_main.ALU_Out_0_4_LC_5_15_5 .LUT_INIT=16'b1000100001100110;
    LogicCell40 \ALU_main.ALU_Out_0_4_LC_5_15_5  (
            .in0(N__7909),
            .in1(N__6209),
            .in2(_gnd_net_),
            .in3(N__6192),
            .lcout(\ALU_main.N_45 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \buf1.out_1_1_iv_LC_5_15_7 .C_ON=1'b0;
    defparam \buf1.out_1_1_iv_LC_5_15_7 .SEQ_MODE=4'b0000;
    defparam \buf1.out_1_1_iv_LC_5_15_7 .LUT_INIT=16'b1111101011111011;
    LogicCell40 \buf1.out_1_1_iv_LC_5_15_7  (
            .in0(N__6635),
            .in1(N__6600),
            .in2(N__6690),
            .in3(N__6551),
            .lcout(bus_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \IR.ff2.q_ner_LC_6_9_1 .C_ON=1'b0;
    defparam \IR.ff2.q_ner_LC_6_9_1 .SEQ_MODE=4'b1010;
    defparam \IR.ff2.q_ner_LC_6_9_1 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \IR.ff2.q_ner_LC_6_9_1  (
            .in0(N__8211),
            .in1(N__8168),
            .in2(N__8121),
            .in3(N__8064),
            .lcout(ir_out_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVIR.ff2.q_nerC_net ),
            .ce(N__8678),
            .sr(N__7297));
    defparam \IR.ff3.q_ner_LC_6_9_2 .C_ON=1'b0;
    defparam \IR.ff3.q_ner_LC_6_9_2 .SEQ_MODE=4'b1010;
    defparam \IR.ff3.q_ner_LC_6_9_2 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \IR.ff3.q_ner_LC_6_9_2  (
            .in0(N__8425),
            .in1(N__8457),
            .in2(N__8368),
            .in3(N__8293),
            .lcout(ir_out_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVIR.ff2.q_nerC_net ),
            .ce(N__8678),
            .sr(N__7297));
    defparam \acc.ff1.q_LC_6_10_0 .C_ON=1'b0;
    defparam \acc.ff1.q_LC_6_10_0 .SEQ_MODE=4'b1010;
    defparam \acc.ff1.q_LC_6_10_0 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \acc.ff1.q_LC_6_10_0  (
            .in0(N__8919),
            .in1(N__8731),
            .in2(N__8860),
            .in3(N__8794),
            .lcout(acc_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVacc.ff1.qC_net ),
            .ce(N__5947),
            .sr(N__7305));
    defparam \acc.ff2.q_LC_6_10_1 .C_ON=1'b0;
    defparam \acc.ff2.q_LC_6_10_1 .SEQ_MODE=4'b1010;
    defparam \acc.ff2.q_LC_6_10_1 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \acc.ff2.q_LC_6_10_1  (
            .in0(N__8167),
            .in1(N__8229),
            .in2(N__8122),
            .in3(N__8053),
            .lcout(acc_out_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVacc.ff1.qC_net ),
            .ce(N__5947),
            .sr(N__7305));
    defparam \acc.ff3.q_LC_6_10_2 .C_ON=1'b0;
    defparam \acc.ff3.q_LC_6_10_2 .SEQ_MODE=4'b1010;
    defparam \acc.ff3.q_LC_6_10_2 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \acc.ff3.q_LC_6_10_2  (
            .in0(N__8306),
            .in1(N__8411),
            .in2(N__8373),
            .in3(N__8478),
            .lcout(acc_out_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVacc.ff1.qC_net ),
            .ce(N__5947),
            .sr(N__7305));
    defparam \acc.ff5.q_LC_6_10_3 .C_ON=1'b0;
    defparam \acc.ff5.q_LC_6_10_3 .SEQ_MODE=4'b1010;
    defparam \acc.ff5.q_LC_6_10_3 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \acc.ff5.q_LC_6_10_3  (
            .in0(N__8003),
            .in1(N__7960),
            .in2(N__7904),
            .in3(N__7479),
            .lcout(acc_out_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVacc.ff1.qC_net ),
            .ce(N__5947),
            .sr(N__7305));
    defparam \mar.ff4.q_ner_LC_6_11_0 .C_ON=1'b0;
    defparam \mar.ff4.q_ner_LC_6_11_0 .SEQ_MODE=4'b1010;
    defparam \mar.ff4.q_ner_LC_6_11_0 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \mar.ff4.q_ner_LC_6_11_0  (
            .in0(N__7748),
            .in1(N__7678),
            .in2(N__7630),
            .in3(N__7546),
            .lcout(mar_out_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVmar.ff4.q_nerC_net ),
            .ce(N__6383),
            .sr(N__7308));
    defparam \mar.ff3.q_ner_LC_6_11_2 .C_ON=1'b0;
    defparam \mar.ff3.q_ner_LC_6_11_2 .SEQ_MODE=4'b1010;
    defparam \mar.ff3.q_ner_LC_6_11_2 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \mar.ff3.q_ner_LC_6_11_2  (
            .in0(N__8426),
            .in1(N__8307),
            .in2(N__8374),
            .in3(N__8479),
            .lcout(mar_out_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVmar.ff4.q_nerC_net ),
            .ce(N__6383),
            .sr(N__7308));
    defparam \mar.ff2.q_ner_LC_6_11_3 .C_ON=1'b0;
    defparam \mar.ff2.q_ner_LC_6_11_3 .SEQ_MODE=4'b1010;
    defparam \mar.ff2.q_ner_LC_6_11_3 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \mar.ff2.q_ner_LC_6_11_3  (
            .in0(N__8236),
            .in1(N__8169),
            .in2(N__8130),
            .in3(N__8052),
            .lcout(mar_out_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVmar.ff4.q_nerC_net ),
            .ce(N__6383),
            .sr(N__7308));
    defparam \b_reg.ff6.q_LC_6_12_0 .C_ON=1'b0;
    defparam \b_reg.ff6.q_LC_6_12_0 .SEQ_MODE=4'b1010;
    defparam \b_reg.ff6.q_LC_6_12_0 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \b_reg.ff6.q_LC_6_12_0  (
            .in0(N__6670),
            .in1(N__6634),
            .in2(N__6598),
            .in3(N__6555),
            .lcout(b_reg_out_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVb_reg.ff6.qC_net ),
            .ce(N__7804),
            .sr(N__7312));
    defparam \b_reg.ff8.q_LC_6_12_1 .C_ON=1'b0;
    defparam \b_reg.ff8.q_LC_6_12_1 .SEQ_MODE=4'b1010;
    defparam \b_reg.ff8.q_LC_6_12_1 .LUT_INIT=16'b1111111111001101;
    LogicCell40 \b_reg.ff8.q_LC_6_12_1  (
            .in0(N__6556),
            .in1(N__6346),
            .in2(N__6890),
            .in3(N__6311),
            .lcout(b_reg_out_7),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVb_reg.ff6.qC_net ),
            .ce(N__7804),
            .sr(N__7312));
    defparam \b_reg.ff1.q_LC_6_12_4 .C_ON=1'b0;
    defparam \b_reg.ff1.q_LC_6_12_4 .SEQ_MODE=4'b1010;
    defparam \b_reg.ff1.q_LC_6_12_4 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \b_reg.ff1.q_LC_6_12_4  (
            .in0(N__8927),
            .in1(N__8848),
            .in2(N__8755),
            .in3(N__8795),
            .lcout(b_reg_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVb_reg.ff6.qC_net ),
            .ce(N__7804),
            .sr(N__7312));
    defparam \mem.data_2_7_0__m18_LC_6_13_0 .C_ON=1'b0;
    defparam \mem.data_2_7_0__m18_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \mem.data_2_7_0__m18_LC_6_13_0 .LUT_INIT=16'b0011111000101111;
    LogicCell40 \mem.data_2_7_0__m18_LC_6_13_0  (
            .in0(N__6962),
            .in1(N__7176),
            .in2(N__7128),
            .in3(N__7029),
            .lcout(),
            .ltout(\mem.i2_mux_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \mem.data_2_7_0__i2_mux_i_m_LC_6_13_1 .C_ON=1'b0;
    defparam \mem.data_2_7_0__i2_mux_i_m_LC_6_13_1 .SEQ_MODE=4'b0000;
    defparam \mem.data_2_7_0__i2_mux_i_m_LC_6_13_1 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \mem.data_2_7_0__i2_mux_i_m_LC_6_13_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6224),
            .in3(N__6553),
            .lcout(mem_data_2_7_0__i2_mux_i_m),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \pc.program_counter_RNO_10_0_LC_6_13_3 .C_ON=1'b0;
    defparam \pc.program_counter_RNO_10_0_LC_6_13_3 .SEQ_MODE=4'b0000;
    defparam \pc.program_counter_RNO_10_0_LC_6_13_3 .LUT_INIT=16'b0111111110011011;
    LogicCell40 \pc.program_counter_RNO_10_0_LC_6_13_3  (
            .in0(N__7175),
            .in1(N__7109),
            .in2(N__7045),
            .in3(N__6960),
            .lcout(\pc.N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \mem.data_2_7_0__m20_LC_6_13_4 .C_ON=1'b0;
    defparam \mem.data_2_7_0__m20_LC_6_13_4 .SEQ_MODE=4'b0000;
    defparam \mem.data_2_7_0__m20_LC_6_13_4 .LUT_INIT=16'b0011111111010111;
    LogicCell40 \mem.data_2_7_0__m20_LC_6_13_4  (
            .in0(N__6961),
            .in1(N__7177),
            .in2(N__7127),
            .in3(N__7028),
            .lcout(m20),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \mem.data_2_7_0__m22_LC_6_13_5 .C_ON=1'b0;
    defparam \mem.data_2_7_0__m22_LC_6_13_5 .SEQ_MODE=4'b0000;
    defparam \mem.data_2_7_0__m22_LC_6_13_5 .LUT_INIT=16'b0111010101110111;
    LogicCell40 \mem.data_2_7_0__m22_LC_6_13_5  (
            .in0(N__7178),
            .in1(N__7114),
            .in2(N__7046),
            .in3(N__6963),
            .lcout(mem_data_2_7_0__N_29_mux),
            .ltout(mem_data_2_7_0__N_29_mux_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \out_reg.ff7.q_LC_6_13_6 .C_ON=1'b0;
    defparam \out_reg.ff7.q_LC_6_13_6 .SEQ_MODE=4'b1010;
    defparam \out_reg.ff7.q_LC_6_13_6 .LUT_INIT=16'b1111111111001101;
    LogicCell40 \out_reg.ff7.q_LC_6_13_6  (
            .in0(N__6554),
            .in1(N__6820),
            .in2(N__7208),
            .in3(N__6782),
            .lcout(out_c_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVout_reg.ff7.qC_net ),
            .ce(N__7473),
            .sr(N__7316));
    defparam \mem.data_2_7_0__m26_LC_6_13_7 .C_ON=1'b0;
    defparam \mem.data_2_7_0__m26_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \mem.data_2_7_0__m26_LC_6_13_7 .LUT_INIT=16'b0001111011111001;
    LogicCell40 \mem.data_2_7_0__m26_LC_6_13_7  (
            .in0(N__7179),
            .in1(N__7113),
            .in2(N__7047),
            .in3(N__6964),
            .lcout(mem_data_2_7_0__i2_mux_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \b_reg.ff2.q_LC_6_14_1 .C_ON=1'b0;
    defparam \b_reg.ff2.q_LC_6_14_1 .SEQ_MODE=4'b1010;
    defparam \b_reg.ff2.q_LC_6_14_1 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \b_reg.ff2.q_LC_6_14_1  (
            .in0(N__8237),
            .in1(N__8183),
            .in2(N__8138),
            .in3(N__8065),
            .lcout(b_reg_out_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVb_reg.ff2.qC_net ),
            .ce(N__7811),
            .sr(N__7320));
    defparam \b_reg.ff7.q_LC_6_14_6 .C_ON=1'b0;
    defparam \b_reg.ff7.q_LC_6_14_6 .SEQ_MODE=4'b1010;
    defparam \b_reg.ff7.q_LC_6_14_6 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \b_reg.ff7.q_LC_6_14_6  (
            .in0(N__6822),
            .in1(N__6790),
            .in2(N__6734),
            .in3(N__6557),
            .lcout(b_reg_out_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVb_reg.ff2.qC_net ),
            .ce(N__7811),
            .sr(N__7320));
    defparam \out_reg.ff6.q_LC_6_15_2 .C_ON=1'b0;
    defparam \out_reg.ff6.q_LC_6_15_2 .SEQ_MODE=4'b1010;
    defparam \out_reg.ff6.q_LC_6_15_2 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \out_reg.ff6.q_LC_6_15_2  (
            .in0(N__6691),
            .in1(N__6637),
            .in2(N__6604),
            .in3(N__6552),
            .lcout(out_c_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVout_reg.ff6.qC_net ),
            .ce(N__7474),
            .sr(N__7322));
    defparam \out_reg.ff3.q_LC_7_9_1 .C_ON=1'b0;
    defparam \out_reg.ff3.q_LC_7_9_1 .SEQ_MODE=4'b1010;
    defparam \out_reg.ff3.q_LC_7_9_1 .LUT_INIT=16'b1111111111001110;
    LogicCell40 \out_reg.ff3.q_LC_7_9_1  (
            .in0(N__8412),
            .in1(N__8468),
            .in2(N__8369),
            .in3(N__8309),
            .lcout(out_c_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVout_reg.ff3.qC_net ),
            .ce(N__7484),
            .sr(N__7302));
    defparam \out_reg.ff1.q_LC_7_9_5 .C_ON=1'b0;
    defparam \out_reg.ff1.q_LC_7_9_5 .SEQ_MODE=4'b1010;
    defparam \out_reg.ff1.q_LC_7_9_5 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \out_reg.ff1.q_LC_7_9_5  (
            .in0(N__8909),
            .in1(N__8732),
            .in2(N__8879),
            .in3(N__8816),
            .lcout(out_c_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVout_reg.ff3.qC_net ),
            .ce(N__7484),
            .sr(N__7302));
    defparam \IR.ff1.q_ner_LC_7_10_0 .C_ON=1'b0;
    defparam \IR.ff1.q_ner_LC_7_10_0 .SEQ_MODE=4'b1010;
    defparam \IR.ff1.q_ner_LC_7_10_0 .LUT_INIT=16'b1111111110111010;
    LogicCell40 \IR.ff1.q_ner_LC_7_10_0  (
            .in0(N__8926),
            .in1(N__8873),
            .in2(N__8748),
            .in3(N__8815),
            .lcout(ir_out_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVIR.ff1.q_nerC_net ),
            .ce(N__8679),
            .sr(N__7309));
    defparam \b_reg.ff3.q_LC_7_11_1 .C_ON=1'b0;
    defparam \b_reg.ff3.q_LC_7_11_1 .SEQ_MODE=4'b1010;
    defparam \b_reg.ff3.q_LC_7_11_1 .LUT_INIT=16'b1111111110101110;
    LogicCell40 \b_reg.ff3.q_LC_7_11_1  (
            .in0(N__8480),
            .in1(N__8427),
            .in2(N__8375),
            .in3(N__8308),
            .lcout(b_reg_out_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVb_reg.ff3.qC_net ),
            .ce(N__7803),
            .sr(N__7313));
    defparam \out_reg.ff2.q_LC_7_12_5 .C_ON=1'b0;
    defparam \out_reg.ff2.q_LC_7_12_5 .SEQ_MODE=4'b1010;
    defparam \out_reg.ff2.q_LC_7_12_5 .LUT_INIT=16'b1111111111011100;
    LogicCell40 \out_reg.ff2.q_LC_7_12_5  (
            .in0(N__8228),
            .in1(N__8182),
            .in2(N__8137),
            .in3(N__8066),
            .lcout(out_c_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVout_reg.ff2.qC_net ),
            .ce(N__7478),
            .sr(N__7317));
    defparam \out_reg.ff5.q_LC_7_12_6 .C_ON=1'b0;
    defparam \out_reg.ff5.q_LC_7_12_6 .SEQ_MODE=4'b1010;
    defparam \out_reg.ff5.q_LC_7_12_6 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \out_reg.ff5.q_LC_7_12_6  (
            .in0(N__8002),
            .in1(N__7952),
            .in2(N__7915),
            .in3(N__7477),
            .lcout(out_c_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVout_reg.ff2.qC_net ),
            .ce(N__7478),
            .sr(N__7317));
    defparam \b_reg.ff4.q_LC_7_13_2 .C_ON=1'b0;
    defparam \b_reg.ff4.q_LC_7_13_2 .SEQ_MODE=4'b1010;
    defparam \b_reg.ff4.q_LC_7_13_2 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \b_reg.ff4.q_LC_7_13_2  (
            .in0(N__7750),
            .in1(N__7685),
            .in2(N__7620),
            .in3(N__7540),
            .lcout(b_reg_out_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVb_reg.ff4.qC_net ),
            .ce(N__7793),
            .sr(N__7321));
    defparam \out_reg.ff4.q_LC_8_11_7 .C_ON=1'b0;
    defparam \out_reg.ff4.q_LC_8_11_7 .SEQ_MODE=4'b1010;
    defparam \out_reg.ff4.q_LC_8_11_7 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \out_reg.ff4.q_LC_8_11_7  (
            .in0(N__7754),
            .in1(N__7679),
            .in2(N__7631),
            .in3(N__7547),
            .lcout(out_c_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVout_reg.ff4.qC_net ),
            .ce(N__7475),
            .sr(N__7318));
endmodule // main
