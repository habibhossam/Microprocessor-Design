-- ******************************************************************************

-- iCEcube Netlister

-- Version:            2020.12.27943

-- Build Date:         Dec  9 2020 18:18:06

-- File Generated:     Dec 13 2023 18:09:27

-- Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

-- Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

-- ******************************************************************************

-- VHDL file for cell "main" view "INTERFACE"

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

library ice;
use ice.vcomponent_vital.all;

-- Entity of main
entity main is
port (
    out : out std_logic_vector(7 downto 0);
    clr : in std_logic;
    clk : in std_logic);
end main;

-- Architecture of main
-- View name is \INTERFACE\
architecture \INTERFACE\ of main is

signal \N__9029\ : std_logic;
signal \N__9028\ : std_logic;
signal \N__9027\ : std_logic;
signal \N__9018\ : std_logic;
signal \N__9017\ : std_logic;
signal \N__9016\ : std_logic;
signal \N__9009\ : std_logic;
signal \N__9008\ : std_logic;
signal \N__9007\ : std_logic;
signal \N__9000\ : std_logic;
signal \N__8999\ : std_logic;
signal \N__8998\ : std_logic;
signal \N__8991\ : std_logic;
signal \N__8990\ : std_logic;
signal \N__8989\ : std_logic;
signal \N__8982\ : std_logic;
signal \N__8981\ : std_logic;
signal \N__8980\ : std_logic;
signal \N__8973\ : std_logic;
signal \N__8972\ : std_logic;
signal \N__8971\ : std_logic;
signal \N__8964\ : std_logic;
signal \N__8963\ : std_logic;
signal \N__8962\ : std_logic;
signal \N__8955\ : std_logic;
signal \N__8954\ : std_logic;
signal \N__8953\ : std_logic;
signal \N__8946\ : std_logic;
signal \N__8945\ : std_logic;
signal \N__8944\ : std_logic;
signal \N__8927\ : std_logic;
signal \N__8926\ : std_logic;
signal \N__8923\ : std_logic;
signal \N__8920\ : std_logic;
signal \N__8919\ : std_logic;
signal \N__8916\ : std_logic;
signal \N__8913\ : std_logic;
signal \N__8910\ : std_logic;
signal \N__8909\ : std_logic;
signal \N__8908\ : std_logic;
signal \N__8901\ : std_logic;
signal \N__8898\ : std_logic;
signal \N__8895\ : std_logic;
signal \N__8892\ : std_logic;
signal \N__8889\ : std_logic;
signal \N__8886\ : std_logic;
signal \N__8879\ : std_logic;
signal \N__8878\ : std_logic;
signal \N__8877\ : std_logic;
signal \N__8874\ : std_logic;
signal \N__8873\ : std_logic;
signal \N__8870\ : std_logic;
signal \N__8867\ : std_logic;
signal \N__8864\ : std_logic;
signal \N__8861\ : std_logic;
signal \N__8860\ : std_logic;
signal \N__8857\ : std_logic;
signal \N__8854\ : std_logic;
signal \N__8849\ : std_logic;
signal \N__8848\ : std_logic;
signal \N__8845\ : std_logic;
signal \N__8842\ : std_logic;
signal \N__8839\ : std_logic;
signal \N__8836\ : std_logic;
signal \N__8833\ : std_logic;
signal \N__8830\ : std_logic;
signal \N__8825\ : std_logic;
signal \N__8816\ : std_logic;
signal \N__8815\ : std_logic;
signal \N__8814\ : std_logic;
signal \N__8811\ : std_logic;
signal \N__8808\ : std_logic;
signal \N__8807\ : std_logic;
signal \N__8804\ : std_logic;
signal \N__8799\ : std_logic;
signal \N__8796\ : std_logic;
signal \N__8795\ : std_logic;
signal \N__8794\ : std_logic;
signal \N__8791\ : std_logic;
signal \N__8788\ : std_logic;
signal \N__8785\ : std_logic;
signal \N__8782\ : std_logic;
signal \N__8779\ : std_logic;
signal \N__8776\ : std_logic;
signal \N__8765\ : std_logic;
signal \N__8764\ : std_logic;
signal \N__8763\ : std_logic;
signal \N__8760\ : std_logic;
signal \N__8757\ : std_logic;
signal \N__8756\ : std_logic;
signal \N__8755\ : std_logic;
signal \N__8752\ : std_logic;
signal \N__8749\ : std_logic;
signal \N__8748\ : std_logic;
signal \N__8745\ : std_logic;
signal \N__8742\ : std_logic;
signal \N__8739\ : std_logic;
signal \N__8736\ : std_logic;
signal \N__8733\ : std_logic;
signal \N__8732\ : std_logic;
signal \N__8731\ : std_logic;
signal \N__8728\ : std_logic;
signal \N__8723\ : std_logic;
signal \N__8720\ : std_logic;
signal \N__8715\ : std_logic;
signal \N__8712\ : std_logic;
signal \N__8709\ : std_logic;
signal \N__8706\ : std_logic;
signal \N__8703\ : std_logic;
signal \N__8698\ : std_logic;
signal \N__8687\ : std_logic;
signal \N__8686\ : std_logic;
signal \N__8685\ : std_logic;
signal \N__8684\ : std_logic;
signal \N__8683\ : std_logic;
signal \N__8680\ : std_logic;
signal \N__8679\ : std_logic;
signal \N__8678\ : std_logic;
signal \N__8677\ : std_logic;
signal \N__8676\ : std_logic;
signal \N__8675\ : std_logic;
signal \N__8674\ : std_logic;
signal \N__8673\ : std_logic;
signal \N__8672\ : std_logic;
signal \N__8669\ : std_logic;
signal \N__8668\ : std_logic;
signal \N__8667\ : std_logic;
signal \N__8666\ : std_logic;
signal \N__8665\ : std_logic;
signal \N__8664\ : std_logic;
signal \N__8663\ : std_logic;
signal \N__8662\ : std_logic;
signal \N__8661\ : std_logic;
signal \N__8660\ : std_logic;
signal \N__8659\ : std_logic;
signal \N__8656\ : std_logic;
signal \N__8655\ : std_logic;
signal \N__8654\ : std_logic;
signal \N__8651\ : std_logic;
signal \N__8648\ : std_logic;
signal \N__8645\ : std_logic;
signal \N__8642\ : std_logic;
signal \N__8639\ : std_logic;
signal \N__8636\ : std_logic;
signal \N__8633\ : std_logic;
signal \N__8630\ : std_logic;
signal \N__8625\ : std_logic;
signal \N__8622\ : std_logic;
signal \N__8621\ : std_logic;
signal \N__8614\ : std_logic;
signal \N__8609\ : std_logic;
signal \N__8604\ : std_logic;
signal \N__8601\ : std_logic;
signal \N__8596\ : std_logic;
signal \N__8587\ : std_logic;
signal \N__8584\ : std_logic;
signal \N__8579\ : std_logic;
signal \N__8576\ : std_logic;
signal \N__8573\ : std_logic;
signal \N__8568\ : std_logic;
signal \N__8563\ : std_logic;
signal \N__8560\ : std_logic;
signal \N__8557\ : std_logic;
signal \N__8554\ : std_logic;
signal \N__8553\ : std_logic;
signal \N__8552\ : std_logic;
signal \N__8551\ : std_logic;
signal \N__8550\ : std_logic;
signal \N__8549\ : std_logic;
signal \N__8548\ : std_logic;
signal \N__8545\ : std_logic;
signal \N__8534\ : std_logic;
signal \N__8531\ : std_logic;
signal \N__8528\ : std_logic;
signal \N__8523\ : std_logic;
signal \N__8514\ : std_logic;
signal \N__8509\ : std_logic;
signal \N__8500\ : std_logic;
signal \N__8495\ : std_logic;
signal \N__8480\ : std_logic;
signal \N__8479\ : std_logic;
signal \N__8478\ : std_logic;
signal \N__8475\ : std_logic;
signal \N__8472\ : std_logic;
signal \N__8469\ : std_logic;
signal \N__8468\ : std_logic;
signal \N__8461\ : std_logic;
signal \N__8458\ : std_logic;
signal \N__8457\ : std_logic;
signal \N__8452\ : std_logic;
signal \N__8449\ : std_logic;
signal \N__8448\ : std_logic;
signal \N__8443\ : std_logic;
signal \N__8440\ : std_logic;
signal \N__8435\ : std_logic;
signal \N__8434\ : std_logic;
signal \N__8431\ : std_logic;
signal \N__8428\ : std_logic;
signal \N__8427\ : std_logic;
signal \N__8426\ : std_logic;
signal \N__8425\ : std_logic;
signal \N__8422\ : std_logic;
signal \N__8419\ : std_logic;
signal \N__8416\ : std_logic;
signal \N__8413\ : std_logic;
signal \N__8412\ : std_logic;
signal \N__8411\ : std_logic;
signal \N__8408\ : std_logic;
signal \N__8403\ : std_logic;
signal \N__8400\ : std_logic;
signal \N__8397\ : std_logic;
signal \N__8394\ : std_logic;
signal \N__8391\ : std_logic;
signal \N__8386\ : std_logic;
signal \N__8375\ : std_logic;
signal \N__8374\ : std_logic;
signal \N__8373\ : std_logic;
signal \N__8370\ : std_logic;
signal \N__8369\ : std_logic;
signal \N__8368\ : std_logic;
signal \N__8365\ : std_logic;
signal \N__8362\ : std_logic;
signal \N__8359\ : std_logic;
signal \N__8356\ : std_logic;
signal \N__8353\ : std_logic;
signal \N__8350\ : std_logic;
signal \N__8347\ : std_logic;
signal \N__8344\ : std_logic;
signal \N__8341\ : std_logic;
signal \N__8338\ : std_logic;
signal \N__8335\ : std_logic;
signal \N__8332\ : std_logic;
signal \N__8325\ : std_logic;
signal \N__8322\ : std_logic;
signal \N__8319\ : std_logic;
signal \N__8316\ : std_logic;
signal \N__8309\ : std_logic;
signal \N__8308\ : std_logic;
signal \N__8307\ : std_logic;
signal \N__8306\ : std_logic;
signal \N__8303\ : std_logic;
signal \N__8300\ : std_logic;
signal \N__8297\ : std_logic;
signal \N__8294\ : std_logic;
signal \N__8293\ : std_logic;
signal \N__8290\ : std_logic;
signal \N__8283\ : std_logic;
signal \N__8280\ : std_logic;
signal \N__8279\ : std_logic;
signal \N__8272\ : std_logic;
signal \N__8269\ : std_logic;
signal \N__8266\ : std_logic;
signal \N__8263\ : std_logic;
signal \N__8258\ : std_logic;
signal \N__8257\ : std_logic;
signal \N__8254\ : std_logic;
signal \N__8253\ : std_logic;
signal \N__8246\ : std_logic;
signal \N__8243\ : std_logic;
signal \N__8240\ : std_logic;
signal \N__8237\ : std_logic;
signal \N__8236\ : std_logic;
signal \N__8233\ : std_logic;
signal \N__8230\ : std_logic;
signal \N__8229\ : std_logic;
signal \N__8228\ : std_logic;
signal \N__8223\ : std_logic;
signal \N__8220\ : std_logic;
signal \N__8217\ : std_logic;
signal \N__8212\ : std_logic;
signal \N__8211\ : std_logic;
signal \N__8210\ : std_logic;
signal \N__8207\ : std_logic;
signal \N__8204\ : std_logic;
signal \N__8201\ : std_logic;
signal \N__8198\ : std_logic;
signal \N__8193\ : std_logic;
signal \N__8188\ : std_logic;
signal \N__8183\ : std_logic;
signal \N__8182\ : std_logic;
signal \N__8179\ : std_logic;
signal \N__8176\ : std_logic;
signal \N__8173\ : std_logic;
signal \N__8170\ : std_logic;
signal \N__8169\ : std_logic;
signal \N__8168\ : std_logic;
signal \N__8167\ : std_logic;
signal \N__8166\ : std_logic;
signal \N__8161\ : std_logic;
signal \N__8158\ : std_logic;
signal \N__8155\ : std_logic;
signal \N__8152\ : std_logic;
signal \N__8149\ : std_logic;
signal \N__8138\ : std_logic;
signal \N__8137\ : std_logic;
signal \N__8134\ : std_logic;
signal \N__8131\ : std_logic;
signal \N__8130\ : std_logic;
signal \N__8129\ : std_logic;
signal \N__8126\ : std_logic;
signal \N__8123\ : std_logic;
signal \N__8122\ : std_logic;
signal \N__8121\ : std_logic;
signal \N__8118\ : std_logic;
signal \N__8115\ : std_logic;
signal \N__8114\ : std_logic;
signal \N__8109\ : std_logic;
signal \N__8106\ : std_logic;
signal \N__8103\ : std_logic;
signal \N__8100\ : std_logic;
signal \N__8097\ : std_logic;
signal \N__8094\ : std_logic;
signal \N__8091\ : std_logic;
signal \N__8088\ : std_logic;
signal \N__8085\ : std_logic;
signal \N__8080\ : std_logic;
signal \N__8077\ : std_logic;
signal \N__8066\ : std_logic;
signal \N__8065\ : std_logic;
signal \N__8064\ : std_logic;
signal \N__8061\ : std_logic;
signal \N__8060\ : std_logic;
signal \N__8057\ : std_logic;
signal \N__8054\ : std_logic;
signal \N__8053\ : std_logic;
signal \N__8052\ : std_logic;
signal \N__8049\ : std_logic;
signal \N__8046\ : std_logic;
signal \N__8045\ : std_logic;
signal \N__8042\ : std_logic;
signal \N__8039\ : std_logic;
signal \N__8036\ : std_logic;
signal \N__8033\ : std_logic;
signal \N__8028\ : std_logic;
signal \N__8025\ : std_logic;
signal \N__8012\ : std_logic;
signal \N__8009\ : std_logic;
signal \N__8006\ : std_logic;
signal \N__8003\ : std_logic;
signal \N__8002\ : std_logic;
signal \N__7999\ : std_logic;
signal \N__7996\ : std_logic;
signal \N__7995\ : std_logic;
signal \N__7994\ : std_logic;
signal \N__7991\ : std_logic;
signal \N__7988\ : std_logic;
signal \N__7985\ : std_logic;
signal \N__7982\ : std_logic;
signal \N__7977\ : std_logic;
signal \N__7974\ : std_logic;
signal \N__7971\ : std_logic;
signal \N__7964\ : std_logic;
signal \N__7961\ : std_logic;
signal \N__7960\ : std_logic;
signal \N__7959\ : std_logic;
signal \N__7956\ : std_logic;
signal \N__7953\ : std_logic;
signal \N__7952\ : std_logic;
signal \N__7951\ : std_logic;
signal \N__7948\ : std_logic;
signal \N__7945\ : std_logic;
signal \N__7942\ : std_logic;
signal \N__7939\ : std_logic;
signal \N__7936\ : std_logic;
signal \N__7933\ : std_logic;
signal \N__7922\ : std_logic;
signal \N__7919\ : std_logic;
signal \N__7916\ : std_logic;
signal \N__7915\ : std_logic;
signal \N__7914\ : std_logic;
signal \N__7911\ : std_logic;
signal \N__7910\ : std_logic;
signal \N__7909\ : std_logic;
signal \N__7908\ : std_logic;
signal \N__7905\ : std_logic;
signal \N__7904\ : std_logic;
signal \N__7903\ : std_logic;
signal \N__7900\ : std_logic;
signal \N__7897\ : std_logic;
signal \N__7892\ : std_logic;
signal \N__7889\ : std_logic;
signal \N__7886\ : std_logic;
signal \N__7883\ : std_logic;
signal \N__7878\ : std_logic;
signal \N__7873\ : std_logic;
signal \N__7870\ : std_logic;
signal \N__7867\ : std_logic;
signal \N__7864\ : std_logic;
signal \N__7857\ : std_logic;
signal \N__7854\ : std_logic;
signal \N__7849\ : std_logic;
signal \N__7844\ : std_logic;
signal \N__7841\ : std_logic;
signal \N__7838\ : std_logic;
signal \N__7835\ : std_logic;
signal \N__7834\ : std_logic;
signal \N__7833\ : std_logic;
signal \N__7830\ : std_logic;
signal \N__7825\ : std_logic;
signal \N__7822\ : std_logic;
signal \N__7819\ : std_logic;
signal \N__7816\ : std_logic;
signal \N__7811\ : std_logic;
signal \N__7808\ : std_logic;
signal \N__7805\ : std_logic;
signal \N__7804\ : std_logic;
signal \N__7803\ : std_logic;
signal \N__7800\ : std_logic;
signal \N__7797\ : std_logic;
signal \N__7794\ : std_logic;
signal \N__7793\ : std_logic;
signal \N__7788\ : std_logic;
signal \N__7785\ : std_logic;
signal \N__7782\ : std_logic;
signal \N__7781\ : std_logic;
signal \N__7778\ : std_logic;
signal \N__7773\ : std_logic;
signal \N__7770\ : std_logic;
signal \N__7767\ : std_logic;
signal \N__7764\ : std_logic;
signal \N__7761\ : std_logic;
signal \N__7754\ : std_logic;
signal \N__7751\ : std_logic;
signal \N__7750\ : std_logic;
signal \N__7749\ : std_logic;
signal \N__7748\ : std_logic;
signal \N__7745\ : std_logic;
signal \N__7742\ : std_logic;
signal \N__7741\ : std_logic;
signal \N__7740\ : std_logic;
signal \N__7737\ : std_logic;
signal \N__7734\ : std_logic;
signal \N__7729\ : std_logic;
signal \N__7726\ : std_logic;
signal \N__7723\ : std_logic;
signal \N__7720\ : std_logic;
signal \N__7717\ : std_logic;
signal \N__7714\ : std_logic;
signal \N__7711\ : std_logic;
signal \N__7706\ : std_logic;
signal \N__7703\ : std_logic;
signal \N__7700\ : std_logic;
signal \N__7697\ : std_logic;
signal \N__7694\ : std_logic;
signal \N__7685\ : std_logic;
signal \N__7682\ : std_logic;
signal \N__7681\ : std_logic;
signal \N__7680\ : std_logic;
signal \N__7679\ : std_logic;
signal \N__7678\ : std_logic;
signal \N__7675\ : std_logic;
signal \N__7672\ : std_logic;
signal \N__7669\ : std_logic;
signal \N__7666\ : std_logic;
signal \N__7663\ : std_logic;
signal \N__7660\ : std_logic;
signal \N__7657\ : std_logic;
signal \N__7654\ : std_logic;
signal \N__7649\ : std_logic;
signal \N__7646\ : std_logic;
signal \N__7643\ : std_logic;
signal \N__7638\ : std_logic;
signal \N__7631\ : std_logic;
signal \N__7630\ : std_logic;
signal \N__7627\ : std_logic;
signal \N__7624\ : std_logic;
signal \N__7621\ : std_logic;
signal \N__7620\ : std_logic;
signal \N__7619\ : std_logic;
signal \N__7618\ : std_logic;
signal \N__7615\ : std_logic;
signal \N__7612\ : std_logic;
signal \N__7609\ : std_logic;
signal \N__7606\ : std_logic;
signal \N__7603\ : std_logic;
signal \N__7600\ : std_logic;
signal \N__7597\ : std_logic;
signal \N__7594\ : std_logic;
signal \N__7593\ : std_logic;
signal \N__7590\ : std_logic;
signal \N__7587\ : std_logic;
signal \N__7584\ : std_logic;
signal \N__7579\ : std_logic;
signal \N__7576\ : std_logic;
signal \N__7573\ : std_logic;
signal \N__7570\ : std_logic;
signal \N__7567\ : std_logic;
signal \N__7564\ : std_logic;
signal \N__7561\ : std_logic;
signal \N__7556\ : std_logic;
signal \N__7547\ : std_logic;
signal \N__7546\ : std_logic;
signal \N__7545\ : std_logic;
signal \N__7544\ : std_logic;
signal \N__7541\ : std_logic;
signal \N__7540\ : std_logic;
signal \N__7537\ : std_logic;
signal \N__7534\ : std_logic;
signal \N__7531\ : std_logic;
signal \N__7528\ : std_logic;
signal \N__7525\ : std_logic;
signal \N__7524\ : std_logic;
signal \N__7521\ : std_logic;
signal \N__7518\ : std_logic;
signal \N__7515\ : std_logic;
signal \N__7510\ : std_logic;
signal \N__7507\ : std_logic;
signal \N__7500\ : std_logic;
signal \N__7493\ : std_logic;
signal \N__7490\ : std_logic;
signal \N__7487\ : std_logic;
signal \N__7484\ : std_logic;
signal \N__7481\ : std_logic;
signal \N__7480\ : std_logic;
signal \N__7479\ : std_logic;
signal \N__7478\ : std_logic;
signal \N__7477\ : std_logic;
signal \N__7476\ : std_logic;
signal \N__7475\ : std_logic;
signal \N__7474\ : std_logic;
signal \N__7473\ : std_logic;
signal \N__7470\ : std_logic;
signal \N__7467\ : std_logic;
signal \N__7464\ : std_logic;
signal \N__7461\ : std_logic;
signal \N__7458\ : std_logic;
signal \N__7457\ : std_logic;
signal \N__7456\ : std_logic;
signal \N__7455\ : std_logic;
signal \N__7454\ : std_logic;
signal \N__7451\ : std_logic;
signal \N__7448\ : std_logic;
signal \N__7445\ : std_logic;
signal \N__7442\ : std_logic;
signal \N__7441\ : std_logic;
signal \N__7438\ : std_logic;
signal \N__7435\ : std_logic;
signal \N__7432\ : std_logic;
signal \N__7427\ : std_logic;
signal \N__7424\ : std_logic;
signal \N__7419\ : std_logic;
signal \N__7416\ : std_logic;
signal \N__7413\ : std_logic;
signal \N__7412\ : std_logic;
signal \N__7409\ : std_logic;
signal \N__7404\ : std_logic;
signal \N__7401\ : std_logic;
signal \N__7400\ : std_logic;
signal \N__7399\ : std_logic;
signal \N__7398\ : std_logic;
signal \N__7389\ : std_logic;
signal \N__7388\ : std_logic;
signal \N__7385\ : std_logic;
signal \N__7378\ : std_logic;
signal \N__7375\ : std_logic;
signal \N__7370\ : std_logic;
signal \N__7367\ : std_logic;
signal \N__7364\ : std_logic;
signal \N__7361\ : std_logic;
signal \N__7358\ : std_logic;
signal \N__7355\ : std_logic;
signal \N__7352\ : std_logic;
signal \N__7345\ : std_logic;
signal \N__7340\ : std_logic;
signal \N__7333\ : std_logic;
signal \N__7322\ : std_logic;
signal \N__7321\ : std_logic;
signal \N__7320\ : std_logic;
signal \N__7319\ : std_logic;
signal \N__7318\ : std_logic;
signal \N__7317\ : std_logic;
signal \N__7316\ : std_logic;
signal \N__7315\ : std_logic;
signal \N__7314\ : std_logic;
signal \N__7313\ : std_logic;
signal \N__7312\ : std_logic;
signal \N__7311\ : std_logic;
signal \N__7310\ : std_logic;
signal \N__7309\ : std_logic;
signal \N__7308\ : std_logic;
signal \N__7307\ : std_logic;
signal \N__7306\ : std_logic;
signal \N__7305\ : std_logic;
signal \N__7304\ : std_logic;
signal \N__7303\ : std_logic;
signal \N__7302\ : std_logic;
signal \N__7301\ : std_logic;
signal \N__7300\ : std_logic;
signal \N__7299\ : std_logic;
signal \N__7298\ : std_logic;
signal \N__7297\ : std_logic;
signal \N__7296\ : std_logic;
signal \N__7295\ : std_logic;
signal \N__7294\ : std_logic;
signal \N__7293\ : std_logic;
signal \N__7292\ : std_logic;
signal \N__7291\ : std_logic;
signal \N__7290\ : std_logic;
signal \N__7289\ : std_logic;
signal \N__7288\ : std_logic;
signal \N__7287\ : std_logic;
signal \N__7214\ : std_logic;
signal \N__7211\ : std_logic;
signal \N__7208\ : std_logic;
signal \N__7205\ : std_logic;
signal \N__7202\ : std_logic;
signal \N__7199\ : std_logic;
signal \N__7196\ : std_logic;
signal \N__7193\ : std_logic;
signal \N__7192\ : std_logic;
signal \N__7187\ : std_logic;
signal \N__7186\ : std_logic;
signal \N__7183\ : std_logic;
signal \N__7180\ : std_logic;
signal \N__7179\ : std_logic;
signal \N__7178\ : std_logic;
signal \N__7177\ : std_logic;
signal \N__7176\ : std_logic;
signal \N__7175\ : std_logic;
signal \N__7174\ : std_logic;
signal \N__7173\ : std_logic;
signal \N__7168\ : std_logic;
signal \N__7167\ : std_logic;
signal \N__7156\ : std_logic;
signal \N__7151\ : std_logic;
signal \N__7148\ : std_logic;
signal \N__7145\ : std_logic;
signal \N__7142\ : std_logic;
signal \N__7139\ : std_logic;
signal \N__7130\ : std_logic;
signal \N__7129\ : std_logic;
signal \N__7128\ : std_logic;
signal \N__7127\ : std_logic;
signal \N__7122\ : std_logic;
signal \N__7121\ : std_logic;
signal \N__7120\ : std_logic;
signal \N__7119\ : std_logic;
signal \N__7118\ : std_logic;
signal \N__7115\ : std_logic;
signal \N__7114\ : std_logic;
signal \N__7113\ : std_logic;
signal \N__7110\ : std_logic;
signal \N__7109\ : std_logic;
signal \N__7108\ : std_logic;
signal \N__7105\ : std_logic;
signal \N__7102\ : std_logic;
signal \N__7099\ : std_logic;
signal \N__7094\ : std_logic;
signal \N__7083\ : std_logic;
signal \N__7080\ : std_logic;
signal \N__7077\ : std_logic;
signal \N__7070\ : std_logic;
signal \N__7067\ : std_logic;
signal \N__7058\ : std_logic;
signal \N__7057\ : std_logic;
signal \N__7054\ : std_logic;
signal \N__7053\ : std_logic;
signal \N__7048\ : std_logic;
signal \N__7047\ : std_logic;
signal \N__7046\ : std_logic;
signal \N__7045\ : std_logic;
signal \N__7044\ : std_logic;
signal \N__7043\ : std_logic;
signal \N__7042\ : std_logic;
signal \N__7039\ : std_logic;
signal \N__7036\ : std_logic;
signal \N__7033\ : std_logic;
signal \N__7030\ : std_logic;
signal \N__7029\ : std_logic;
signal \N__7028\ : std_logic;
signal \N__7025\ : std_logic;
signal \N__7022\ : std_logic;
signal \N__7019\ : std_logic;
signal \N__7018\ : std_logic;
signal \N__7015\ : std_logic;
signal \N__7012\ : std_logic;
signal \N__7009\ : std_logic;
signal \N__6998\ : std_logic;
signal \N__6995\ : std_logic;
signal \N__6988\ : std_logic;
signal \N__6985\ : std_logic;
signal \N__6980\ : std_logic;
signal \N__6975\ : std_logic;
signal \N__6968\ : std_logic;
signal \N__6967\ : std_logic;
signal \N__6966\ : std_logic;
signal \N__6965\ : std_logic;
signal \N__6964\ : std_logic;
signal \N__6963\ : std_logic;
signal \N__6962\ : std_logic;
signal \N__6961\ : std_logic;
signal \N__6960\ : std_logic;
signal \N__6957\ : std_logic;
signal \N__6952\ : std_logic;
signal \N__6949\ : std_logic;
signal \N__6938\ : std_logic;
signal \N__6935\ : std_logic;
signal \N__6934\ : std_logic;
signal \N__6933\ : std_logic;
signal \N__6932\ : std_logic;
signal \N__6927\ : std_logic;
signal \N__6924\ : std_logic;
signal \N__6921\ : std_logic;
signal \N__6914\ : std_logic;
signal \N__6909\ : std_logic;
signal \N__6902\ : std_logic;
signal \N__6901\ : std_logic;
signal \N__6900\ : std_logic;
signal \N__6895\ : std_logic;
signal \N__6892\ : std_logic;
signal \N__6891\ : std_logic;
signal \N__6890\ : std_logic;
signal \N__6887\ : std_logic;
signal \N__6884\ : std_logic;
signal \N__6881\ : std_logic;
signal \N__6878\ : std_logic;
signal \N__6875\ : std_logic;
signal \N__6872\ : std_logic;
signal \N__6869\ : std_logic;
signal \N__6866\ : std_logic;
signal \N__6863\ : std_logic;
signal \N__6854\ : std_logic;
signal \N__6851\ : std_logic;
signal \N__6848\ : std_logic;
signal \N__6847\ : std_logic;
signal \N__6844\ : std_logic;
signal \N__6841\ : std_logic;
signal \N__6836\ : std_logic;
signal \N__6833\ : std_logic;
signal \N__6830\ : std_logic;
signal \N__6829\ : std_logic;
signal \N__6826\ : std_logic;
signal \N__6823\ : std_logic;
signal \N__6822\ : std_logic;
signal \N__6821\ : std_logic;
signal \N__6820\ : std_logic;
signal \N__6817\ : std_logic;
signal \N__6814\ : std_logic;
signal \N__6811\ : std_logic;
signal \N__6808\ : std_logic;
signal \N__6805\ : std_logic;
signal \N__6800\ : std_logic;
signal \N__6791\ : std_logic;
signal \N__6790\ : std_logic;
signal \N__6789\ : std_logic;
signal \N__6786\ : std_logic;
signal \N__6783\ : std_logic;
signal \N__6782\ : std_logic;
signal \N__6779\ : std_logic;
signal \N__6778\ : std_logic;
signal \N__6775\ : std_logic;
signal \N__6772\ : std_logic;
signal \N__6769\ : std_logic;
signal \N__6766\ : std_logic;
signal \N__6763\ : std_logic;
signal \N__6756\ : std_logic;
signal \N__6753\ : std_logic;
signal \N__6746\ : std_logic;
signal \N__6745\ : std_logic;
signal \N__6742\ : std_logic;
signal \N__6739\ : std_logic;
signal \N__6736\ : std_logic;
signal \N__6735\ : std_logic;
signal \N__6734\ : std_logic;
signal \N__6729\ : std_logic;
signal \N__6726\ : std_logic;
signal \N__6723\ : std_logic;
signal \N__6720\ : std_logic;
signal \N__6717\ : std_logic;
signal \N__6714\ : std_logic;
signal \N__6711\ : std_logic;
signal \N__6704\ : std_logic;
signal \N__6703\ : std_logic;
signal \N__6700\ : std_logic;
signal \N__6697\ : std_logic;
signal \N__6692\ : std_logic;
signal \N__6691\ : std_logic;
signal \N__6690\ : std_logic;
signal \N__6687\ : std_logic;
signal \N__6684\ : std_logic;
signal \N__6683\ : std_logic;
signal \N__6680\ : std_logic;
signal \N__6677\ : std_logic;
signal \N__6674\ : std_logic;
signal \N__6671\ : std_logic;
signal \N__6670\ : std_logic;
signal \N__6667\ : std_logic;
signal \N__6664\ : std_logic;
signal \N__6661\ : std_logic;
signal \N__6658\ : std_logic;
signal \N__6655\ : std_logic;
signal \N__6652\ : std_logic;
signal \N__6641\ : std_logic;
signal \N__6638\ : std_logic;
signal \N__6637\ : std_logic;
signal \N__6636\ : std_logic;
signal \N__6635\ : std_logic;
signal \N__6634\ : std_logic;
signal \N__6631\ : std_logic;
signal \N__6628\ : std_logic;
signal \N__6625\ : std_logic;
signal \N__6622\ : std_logic;
signal \N__6619\ : std_logic;
signal \N__6610\ : std_logic;
signal \N__6605\ : std_logic;
signal \N__6604\ : std_logic;
signal \N__6601\ : std_logic;
signal \N__6600\ : std_logic;
signal \N__6599\ : std_logic;
signal \N__6598\ : std_logic;
signal \N__6595\ : std_logic;
signal \N__6592\ : std_logic;
signal \N__6589\ : std_logic;
signal \N__6586\ : std_logic;
signal \N__6583\ : std_logic;
signal \N__6580\ : std_logic;
signal \N__6575\ : std_logic;
signal \N__6572\ : std_logic;
signal \N__6569\ : std_logic;
signal \N__6564\ : std_logic;
signal \N__6557\ : std_logic;
signal \N__6556\ : std_logic;
signal \N__6555\ : std_logic;
signal \N__6554\ : std_logic;
signal \N__6553\ : std_logic;
signal \N__6552\ : std_logic;
signal \N__6551\ : std_logic;
signal \N__6548\ : std_logic;
signal \N__6543\ : std_logic;
signal \N__6538\ : std_logic;
signal \N__6537\ : std_logic;
signal \N__6536\ : std_logic;
signal \N__6535\ : std_logic;
signal \N__6534\ : std_logic;
signal \N__6531\ : std_logic;
signal \N__6528\ : std_logic;
signal \N__6527\ : std_logic;
signal \N__6526\ : std_logic;
signal \N__6525\ : std_logic;
signal \N__6524\ : std_logic;
signal \N__6523\ : std_logic;
signal \N__6522\ : std_logic;
signal \N__6521\ : std_logic;
signal \N__6514\ : std_logic;
signal \N__6511\ : std_logic;
signal \N__6504\ : std_logic;
signal \N__6499\ : std_logic;
signal \N__6496\ : std_logic;
signal \N__6489\ : std_logic;
signal \N__6486\ : std_logic;
signal \N__6483\ : std_logic;
signal \N__6482\ : std_logic;
signal \N__6479\ : std_logic;
signal \N__6474\ : std_logic;
signal \N__6467\ : std_logic;
signal \N__6466\ : std_logic;
signal \N__6465\ : std_logic;
signal \N__6464\ : std_logic;
signal \N__6463\ : std_logic;
signal \N__6460\ : std_logic;
signal \N__6455\ : std_logic;
signal \N__6452\ : std_logic;
signal \N__6445\ : std_logic;
signal \N__6438\ : std_logic;
signal \N__6435\ : std_logic;
signal \N__6422\ : std_logic;
signal \N__6419\ : std_logic;
signal \N__6416\ : std_logic;
signal \N__6413\ : std_logic;
signal \N__6410\ : std_logic;
signal \N__6407\ : std_logic;
signal \N__6404\ : std_logic;
signal \N__6401\ : std_logic;
signal \N__6398\ : std_logic;
signal \N__6395\ : std_logic;
signal \N__6392\ : std_logic;
signal \N__6389\ : std_logic;
signal \N__6386\ : std_logic;
signal \N__6383\ : std_logic;
signal \N__6382\ : std_logic;
signal \N__6379\ : std_logic;
signal \N__6376\ : std_logic;
signal \N__6373\ : std_logic;
signal \N__6370\ : std_logic;
signal \N__6365\ : std_logic;
signal \N__6362\ : std_logic;
signal \N__6359\ : std_logic;
signal \N__6358\ : std_logic;
signal \N__6353\ : std_logic;
signal \N__6350\ : std_logic;
signal \N__6347\ : std_logic;
signal \N__6346\ : std_logic;
signal \N__6343\ : std_logic;
signal \N__6340\ : std_logic;
signal \N__6335\ : std_logic;
signal \N__6334\ : std_logic;
signal \N__6331\ : std_logic;
signal \N__6328\ : std_logic;
signal \N__6327\ : std_logic;
signal \N__6324\ : std_logic;
signal \N__6321\ : std_logic;
signal \N__6318\ : std_logic;
signal \N__6311\ : std_logic;
signal \N__6310\ : std_logic;
signal \N__6309\ : std_logic;
signal \N__6306\ : std_logic;
signal \N__6303\ : std_logic;
signal \N__6300\ : std_logic;
signal \N__6297\ : std_logic;
signal \N__6294\ : std_logic;
signal \N__6293\ : std_logic;
signal \N__6290\ : std_logic;
signal \N__6285\ : std_logic;
signal \N__6282\ : std_logic;
signal \N__6279\ : std_logic;
signal \N__6276\ : std_logic;
signal \N__6269\ : std_logic;
signal \N__6268\ : std_logic;
signal \N__6265\ : std_logic;
signal \N__6262\ : std_logic;
signal \N__6259\ : std_logic;
signal \N__6256\ : std_logic;
signal \N__6251\ : std_logic;
signal \N__6248\ : std_logic;
signal \N__6245\ : std_logic;
signal \N__6244\ : std_logic;
signal \N__6243\ : std_logic;
signal \N__6240\ : std_logic;
signal \N__6235\ : std_logic;
signal \N__6232\ : std_logic;
signal \N__6229\ : std_logic;
signal \N__6224\ : std_logic;
signal \N__6221\ : std_logic;
signal \N__6218\ : std_logic;
signal \N__6215\ : std_logic;
signal \N__6212\ : std_logic;
signal \N__6209\ : std_logic;
signal \N__6206\ : std_logic;
signal \N__6205\ : std_logic;
signal \N__6202\ : std_logic;
signal \N__6199\ : std_logic;
signal \N__6194\ : std_logic;
signal \N__6193\ : std_logic;
signal \N__6192\ : std_logic;
signal \N__6191\ : std_logic;
signal \N__6190\ : std_logic;
signal \N__6187\ : std_logic;
signal \N__6186\ : std_logic;
signal \N__6183\ : std_logic;
signal \N__6180\ : std_logic;
signal \N__6175\ : std_logic;
signal \N__6172\ : std_logic;
signal \N__6169\ : std_logic;
signal \N__6168\ : std_logic;
signal \N__6167\ : std_logic;
signal \N__6166\ : std_logic;
signal \N__6165\ : std_logic;
signal \N__6164\ : std_logic;
signal \N__6163\ : std_logic;
signal \N__6162\ : std_logic;
signal \N__6161\ : std_logic;
signal \N__6160\ : std_logic;
signal \N__6159\ : std_logic;
signal \N__6158\ : std_logic;
signal \N__6157\ : std_logic;
signal \N__6156\ : std_logic;
signal \N__6153\ : std_logic;
signal \N__6148\ : std_logic;
signal \N__6143\ : std_logic;
signal \N__6136\ : std_logic;
signal \N__6131\ : std_logic;
signal \N__6124\ : std_logic;
signal \N__6119\ : std_logic;
signal \N__6112\ : std_logic;
signal \N__6095\ : std_logic;
signal \N__6092\ : std_logic;
signal \N__6089\ : std_logic;
signal \N__6086\ : std_logic;
signal \N__6083\ : std_logic;
signal \N__6080\ : std_logic;
signal \N__6079\ : std_logic;
signal \N__6076\ : std_logic;
signal \N__6073\ : std_logic;
signal \N__6068\ : std_logic;
signal \N__6067\ : std_logic;
signal \N__6064\ : std_logic;
signal \N__6061\ : std_logic;
signal \N__6060\ : std_logic;
signal \N__6055\ : std_logic;
signal \N__6052\ : std_logic;
signal \N__6051\ : std_logic;
signal \N__6050\ : std_logic;
signal \N__6045\ : std_logic;
signal \N__6042\ : std_logic;
signal \N__6039\ : std_logic;
signal \N__6036\ : std_logic;
signal \N__6029\ : std_logic;
signal \N__6028\ : std_logic;
signal \N__6025\ : std_logic;
signal \N__6024\ : std_logic;
signal \N__6021\ : std_logic;
signal \N__6018\ : std_logic;
signal \N__6015\ : std_logic;
signal \N__6014\ : std_logic;
signal \N__6011\ : std_logic;
signal \N__6006\ : std_logic;
signal \N__6003\ : std_logic;
signal \N__6000\ : std_logic;
signal \N__5993\ : std_logic;
signal \N__5992\ : std_logic;
signal \N__5991\ : std_logic;
signal \N__5990\ : std_logic;
signal \N__5989\ : std_logic;
signal \N__5986\ : std_logic;
signal \N__5979\ : std_logic;
signal \N__5976\ : std_logic;
signal \N__5973\ : std_logic;
signal \N__5970\ : std_logic;
signal \N__5967\ : std_logic;
signal \N__5964\ : std_logic;
signal \N__5961\ : std_logic;
signal \N__5958\ : std_logic;
signal \N__5955\ : std_logic;
signal \N__5948\ : std_logic;
signal \N__5947\ : std_logic;
signal \N__5944\ : std_logic;
signal \N__5941\ : std_logic;
signal \N__5938\ : std_logic;
signal \N__5935\ : std_logic;
signal \N__5932\ : std_logic;
signal \N__5929\ : std_logic;
signal \N__5924\ : std_logic;
signal \N__5921\ : std_logic;
signal \N__5918\ : std_logic;
signal \N__5915\ : std_logic;
signal \N__5912\ : std_logic;
signal \N__5909\ : std_logic;
signal \N__5908\ : std_logic;
signal \N__5907\ : std_logic;
signal \N__5906\ : std_logic;
signal \N__5903\ : std_logic;
signal \N__5900\ : std_logic;
signal \N__5895\ : std_logic;
signal \N__5892\ : std_logic;
signal \N__5885\ : std_logic;
signal \N__5882\ : std_logic;
signal \N__5879\ : std_logic;
signal \N__5876\ : std_logic;
signal \N__5875\ : std_logic;
signal \N__5870\ : std_logic;
signal \N__5867\ : std_logic;
signal \N__5866\ : std_logic;
signal \N__5863\ : std_logic;
signal \N__5860\ : std_logic;
signal \N__5855\ : std_logic;
signal \N__5854\ : std_logic;
signal \N__5853\ : std_logic;
signal \N__5852\ : std_logic;
signal \N__5849\ : std_logic;
signal \N__5842\ : std_logic;
signal \N__5839\ : std_logic;
signal \N__5834\ : std_logic;
signal \N__5831\ : std_logic;
signal \N__5828\ : std_logic;
signal \N__5827\ : std_logic;
signal \N__5824\ : std_logic;
signal \N__5823\ : std_logic;
signal \N__5822\ : std_logic;
signal \N__5821\ : std_logic;
signal \N__5820\ : std_logic;
signal \N__5817\ : std_logic;
signal \N__5814\ : std_logic;
signal \N__5811\ : std_logic;
signal \N__5808\ : std_logic;
signal \N__5803\ : std_logic;
signal \N__5800\ : std_logic;
signal \N__5797\ : std_logic;
signal \N__5794\ : std_logic;
signal \N__5789\ : std_logic;
signal \N__5784\ : std_logic;
signal \N__5777\ : std_logic;
signal \N__5774\ : std_logic;
signal \N__5771\ : std_logic;
signal \N__5768\ : std_logic;
signal \N__5767\ : std_logic;
signal \N__5764\ : std_logic;
signal \N__5763\ : std_logic;
signal \N__5762\ : std_logic;
signal \N__5761\ : std_logic;
signal \N__5760\ : std_logic;
signal \N__5757\ : std_logic;
signal \N__5754\ : std_logic;
signal \N__5749\ : std_logic;
signal \N__5748\ : std_logic;
signal \N__5747\ : std_logic;
signal \N__5746\ : std_logic;
signal \N__5743\ : std_logic;
signal \N__5742\ : std_logic;
signal \N__5741\ : std_logic;
signal \N__5738\ : std_logic;
signal \N__5735\ : std_logic;
signal \N__5732\ : std_logic;
signal \N__5729\ : std_logic;
signal \N__5722\ : std_logic;
signal \N__5719\ : std_logic;
signal \N__5714\ : std_logic;
signal \N__5711\ : std_logic;
signal \N__5702\ : std_logic;
signal \N__5697\ : std_logic;
signal \N__5694\ : std_logic;
signal \N__5689\ : std_logic;
signal \N__5684\ : std_logic;
signal \N__5683\ : std_logic;
signal \N__5682\ : std_logic;
signal \N__5681\ : std_logic;
signal \N__5680\ : std_logic;
signal \N__5679\ : std_logic;
signal \N__5676\ : std_logic;
signal \N__5675\ : std_logic;
signal \N__5674\ : std_logic;
signal \N__5673\ : std_logic;
signal \N__5668\ : std_logic;
signal \N__5665\ : std_logic;
signal \N__5662\ : std_logic;
signal \N__5659\ : std_logic;
signal \N__5656\ : std_logic;
signal \N__5653\ : std_logic;
signal \N__5648\ : std_logic;
signal \N__5645\ : std_logic;
signal \N__5644\ : std_logic;
signal \N__5643\ : std_logic;
signal \N__5640\ : std_logic;
signal \N__5637\ : std_logic;
signal \N__5634\ : std_logic;
signal \N__5631\ : std_logic;
signal \N__5626\ : std_logic;
signal \N__5623\ : std_logic;
signal \N__5618\ : std_logic;
signal \N__5611\ : std_logic;
signal \N__5602\ : std_logic;
signal \N__5597\ : std_logic;
signal \N__5594\ : std_logic;
signal \N__5591\ : std_logic;
signal \N__5590\ : std_logic;
signal \N__5587\ : std_logic;
signal \N__5584\ : std_logic;
signal \N__5581\ : std_logic;
signal \N__5578\ : std_logic;
signal \N__5575\ : std_logic;
signal \N__5572\ : std_logic;
signal \N__5567\ : std_logic;
signal \N__5564\ : std_logic;
signal \N__5563\ : std_logic;
signal \N__5562\ : std_logic;
signal \N__5561\ : std_logic;
signal \N__5558\ : std_logic;
signal \N__5555\ : std_logic;
signal \N__5550\ : std_logic;
signal \N__5549\ : std_logic;
signal \N__5548\ : std_logic;
signal \N__5547\ : std_logic;
signal \N__5546\ : std_logic;
signal \N__5545\ : std_logic;
signal \N__5542\ : std_logic;
signal \N__5539\ : std_logic;
signal \N__5536\ : std_logic;
signal \N__5531\ : std_logic;
signal \N__5526\ : std_logic;
signal \N__5523\ : std_logic;
signal \N__5510\ : std_logic;
signal \N__5507\ : std_logic;
signal \N__5504\ : std_logic;
signal \N__5501\ : std_logic;
signal \N__5500\ : std_logic;
signal \N__5499\ : std_logic;
signal \N__5498\ : std_logic;
signal \N__5497\ : std_logic;
signal \N__5496\ : std_logic;
signal \N__5495\ : std_logic;
signal \N__5494\ : std_logic;
signal \N__5491\ : std_logic;
signal \N__5488\ : std_logic;
signal \N__5483\ : std_logic;
signal \N__5478\ : std_logic;
signal \N__5475\ : std_logic;
signal \N__5472\ : std_logic;
signal \N__5469\ : std_logic;
signal \N__5456\ : std_logic;
signal \N__5455\ : std_logic;
signal \N__5452\ : std_logic;
signal \N__5449\ : std_logic;
signal \N__5448\ : std_logic;
signal \N__5447\ : std_logic;
signal \N__5446\ : std_logic;
signal \N__5445\ : std_logic;
signal \N__5444\ : std_logic;
signal \N__5443\ : std_logic;
signal \N__5440\ : std_logic;
signal \N__5437\ : std_logic;
signal \N__5430\ : std_logic;
signal \N__5427\ : std_logic;
signal \N__5422\ : std_logic;
signal \N__5419\ : std_logic;
signal \N__5408\ : std_logic;
signal \N__5407\ : std_logic;
signal \N__5406\ : std_logic;
signal \N__5405\ : std_logic;
signal \N__5402\ : std_logic;
signal \N__5399\ : std_logic;
signal \N__5398\ : std_logic;
signal \N__5397\ : std_logic;
signal \N__5394\ : std_logic;
signal \N__5391\ : std_logic;
signal \N__5388\ : std_logic;
signal \N__5385\ : std_logic;
signal \N__5380\ : std_logic;
signal \N__5377\ : std_logic;
signal \N__5366\ : std_logic;
signal \N__5365\ : std_logic;
signal \N__5364\ : std_logic;
signal \N__5363\ : std_logic;
signal \N__5362\ : std_logic;
signal \N__5359\ : std_logic;
signal \N__5354\ : std_logic;
signal \N__5351\ : std_logic;
signal \N__5350\ : std_logic;
signal \N__5347\ : std_logic;
signal \N__5342\ : std_logic;
signal \N__5339\ : std_logic;
signal \N__5334\ : std_logic;
signal \N__5327\ : std_logic;
signal \N__5326\ : std_logic;
signal \N__5325\ : std_logic;
signal \N__5322\ : std_logic;
signal \N__5317\ : std_logic;
signal \N__5312\ : std_logic;
signal \N__5311\ : std_logic;
signal \N__5310\ : std_logic;
signal \N__5309\ : std_logic;
signal \N__5306\ : std_logic;
signal \N__5303\ : std_logic;
signal \N__5300\ : std_logic;
signal \N__5299\ : std_logic;
signal \N__5296\ : std_logic;
signal \N__5295\ : std_logic;
signal \N__5292\ : std_logic;
signal \N__5291\ : std_logic;
signal \N__5290\ : std_logic;
signal \N__5285\ : std_logic;
signal \N__5282\ : std_logic;
signal \N__5281\ : std_logic;
signal \N__5278\ : std_logic;
signal \N__5275\ : std_logic;
signal \N__5272\ : std_logic;
signal \N__5267\ : std_logic;
signal \N__5264\ : std_logic;
signal \N__5259\ : std_logic;
signal \N__5246\ : std_logic;
signal \N__5243\ : std_logic;
signal \N__5240\ : std_logic;
signal \N__5237\ : std_logic;
signal \N__5234\ : std_logic;
signal \N__5231\ : std_logic;
signal \N__5228\ : std_logic;
signal \N__5225\ : std_logic;
signal \N__5222\ : std_logic;
signal \N__5219\ : std_logic;
signal \N__5218\ : std_logic;
signal \N__5217\ : std_logic;
signal \N__5216\ : std_logic;
signal \N__5213\ : std_logic;
signal \N__5210\ : std_logic;
signal \N__5207\ : std_logic;
signal \N__5204\ : std_logic;
signal \N__5203\ : std_logic;
signal \N__5202\ : std_logic;
signal \N__5197\ : std_logic;
signal \N__5192\ : std_logic;
signal \N__5189\ : std_logic;
signal \N__5188\ : std_logic;
signal \N__5185\ : std_logic;
signal \N__5182\ : std_logic;
signal \N__5179\ : std_logic;
signal \N__5176\ : std_logic;
signal \N__5173\ : std_logic;
signal \N__5170\ : std_logic;
signal \N__5165\ : std_logic;
signal \N__5156\ : std_logic;
signal \N__5155\ : std_logic;
signal \N__5154\ : std_logic;
signal \N__5151\ : std_logic;
signal \N__5148\ : std_logic;
signal \N__5147\ : std_logic;
signal \N__5144\ : std_logic;
signal \N__5139\ : std_logic;
signal \N__5138\ : std_logic;
signal \N__5135\ : std_logic;
signal \N__5134\ : std_logic;
signal \N__5133\ : std_logic;
signal \N__5130\ : std_logic;
signal \N__5127\ : std_logic;
signal \N__5120\ : std_logic;
signal \N__5117\ : std_logic;
signal \N__5108\ : std_logic;
signal \N__5105\ : std_logic;
signal \N__5102\ : std_logic;
signal \N__5099\ : std_logic;
signal \N__5096\ : std_logic;
signal \N__5093\ : std_logic;
signal \N__5092\ : std_logic;
signal \N__5089\ : std_logic;
signal \N__5088\ : std_logic;
signal \N__5085\ : std_logic;
signal \N__5082\ : std_logic;
signal \N__5079\ : std_logic;
signal \N__5078\ : std_logic;
signal \N__5075\ : std_logic;
signal \N__5070\ : std_logic;
signal \N__5067\ : std_logic;
signal \N__5060\ : std_logic;
signal \N__5057\ : std_logic;
signal \N__5054\ : std_logic;
signal \N__5051\ : std_logic;
signal \N__5048\ : std_logic;
signal \N__5045\ : std_logic;
signal \N__5042\ : std_logic;
signal \N__5039\ : std_logic;
signal \N__5036\ : std_logic;
signal \N__5033\ : std_logic;
signal \N__5030\ : std_logic;
signal \N__5029\ : std_logic;
signal \N__5026\ : std_logic;
signal \N__5023\ : std_logic;
signal \N__5020\ : std_logic;
signal \N__5015\ : std_logic;
signal \N__5014\ : std_logic;
signal \N__5009\ : std_logic;
signal \N__5006\ : std_logic;
signal \N__5005\ : std_logic;
signal \N__5004\ : std_logic;
signal \N__5003\ : std_logic;
signal \N__5002\ : std_logic;
signal \N__4999\ : std_logic;
signal \N__4992\ : std_logic;
signal \N__4989\ : std_logic;
signal \N__4982\ : std_logic;
signal \N__4981\ : std_logic;
signal \N__4980\ : std_logic;
signal \N__4977\ : std_logic;
signal \N__4972\ : std_logic;
signal \N__4969\ : std_logic;
signal \N__4966\ : std_logic;
signal \N__4965\ : std_logic;
signal \N__4964\ : std_logic;
signal \N__4963\ : std_logic;
signal \N__4958\ : std_logic;
signal \N__4953\ : std_logic;
signal \N__4950\ : std_logic;
signal \N__4943\ : std_logic;
signal \N__4940\ : std_logic;
signal \N__4937\ : std_logic;
signal \N__4934\ : std_logic;
signal \N__4931\ : std_logic;
signal \N__4928\ : std_logic;
signal \N__4925\ : std_logic;
signal \N__4922\ : std_logic;
signal \N__4919\ : std_logic;
signal \N__4916\ : std_logic;
signal \N__4913\ : std_logic;
signal \N__4910\ : std_logic;
signal \N__4907\ : std_logic;
signal \N__4904\ : std_logic;
signal \N__4901\ : std_logic;
signal \N__4898\ : std_logic;
signal \N__4897\ : std_logic;
signal \N__4894\ : std_logic;
signal \N__4891\ : std_logic;
signal \N__4890\ : std_logic;
signal \N__4889\ : std_logic;
signal \N__4884\ : std_logic;
signal \N__4879\ : std_logic;
signal \N__4874\ : std_logic;
signal \N__4871\ : std_logic;
signal \N__4868\ : std_logic;
signal \N__4865\ : std_logic;
signal \N__4862\ : std_logic;
signal \N__4859\ : std_logic;
signal \N__4856\ : std_logic;
signal \N__4853\ : std_logic;
signal \N__4850\ : std_logic;
signal \N__4847\ : std_logic;
signal \N__4844\ : std_logic;
signal \N__4841\ : std_logic;
signal \N__4838\ : std_logic;
signal \N__4837\ : std_logic;
signal \N__4834\ : std_logic;
signal \N__4833\ : std_logic;
signal \N__4832\ : std_logic;
signal \N__4829\ : std_logic;
signal \N__4826\ : std_logic;
signal \N__4823\ : std_logic;
signal \N__4820\ : std_logic;
signal \N__4817\ : std_logic;
signal \N__4808\ : std_logic;
signal \N__4807\ : std_logic;
signal \N__4806\ : std_logic;
signal \N__4805\ : std_logic;
signal \N__4804\ : std_logic;
signal \N__4803\ : std_logic;
signal \N__4802\ : std_logic;
signal \N__4801\ : std_logic;
signal \N__4800\ : std_logic;
signal \N__4799\ : std_logic;
signal \N__4798\ : std_logic;
signal \N__4797\ : std_logic;
signal \N__4796\ : std_logic;
signal \N__4795\ : std_logic;
signal \N__4794\ : std_logic;
signal \N__4793\ : std_logic;
signal \N__4792\ : std_logic;
signal \N__4791\ : std_logic;
signal \N__4790\ : std_logic;
signal \N__4789\ : std_logic;
signal \N__4788\ : std_logic;
signal \N__4787\ : std_logic;
signal \N__4786\ : std_logic;
signal \N__4785\ : std_logic;
signal \N__4784\ : std_logic;
signal \N__4783\ : std_logic;
signal \N__4782\ : std_logic;
signal \N__4781\ : std_logic;
signal \N__4780\ : std_logic;
signal \N__4779\ : std_logic;
signal \N__4778\ : std_logic;
signal \N__4777\ : std_logic;
signal \N__4776\ : std_logic;
signal \N__4775\ : std_logic;
signal \N__4774\ : std_logic;
signal \N__4773\ : std_logic;
signal \N__4700\ : std_logic;
signal \N__4697\ : std_logic;
signal \N__4694\ : std_logic;
signal \N__4693\ : std_logic;
signal \N__4692\ : std_logic;
signal \N__4691\ : std_logic;
signal \N__4690\ : std_logic;
signal \N__4687\ : std_logic;
signal \N__4686\ : std_logic;
signal \N__4681\ : std_logic;
signal \N__4678\ : std_logic;
signal \N__4673\ : std_logic;
signal \N__4670\ : std_logic;
signal \N__4669\ : std_logic;
signal \N__4668\ : std_logic;
signal \N__4667\ : std_logic;
signal \N__4666\ : std_logic;
signal \N__4663\ : std_logic;
signal \N__4658\ : std_logic;
signal \N__4655\ : std_logic;
signal \N__4654\ : std_logic;
signal \N__4651\ : std_logic;
signal \N__4648\ : std_logic;
signal \N__4645\ : std_logic;
signal \N__4644\ : std_logic;
signal \N__4641\ : std_logic;
signal \N__4640\ : std_logic;
signal \N__4639\ : std_logic;
signal \N__4632\ : std_logic;
signal \N__4629\ : std_logic;
signal \N__4626\ : std_logic;
signal \N__4623\ : std_logic;
signal \N__4620\ : std_logic;
signal \N__4615\ : std_logic;
signal \N__4610\ : std_logic;
signal \N__4607\ : std_logic;
signal \N__4604\ : std_logic;
signal \N__4589\ : std_logic;
signal \N__4588\ : std_logic;
signal \N__4587\ : std_logic;
signal \N__4584\ : std_logic;
signal \N__4581\ : std_logic;
signal \N__4580\ : std_logic;
signal \N__4579\ : std_logic;
signal \N__4578\ : std_logic;
signal \N__4577\ : std_logic;
signal \N__4574\ : std_logic;
signal \N__4571\ : std_logic;
signal \N__4568\ : std_logic;
signal \N__4563\ : std_logic;
signal \N__4558\ : std_logic;
signal \N__4555\ : std_logic;
signal \N__4548\ : std_logic;
signal \N__4547\ : std_logic;
signal \N__4544\ : std_logic;
signal \N__4543\ : std_logic;
signal \N__4542\ : std_logic;
signal \N__4541\ : std_logic;
signal \N__4540\ : std_logic;
signal \N__4539\ : std_logic;
signal \N__4536\ : std_logic;
signal \N__4533\ : std_logic;
signal \N__4530\ : std_logic;
signal \N__4527\ : std_logic;
signal \N__4522\ : std_logic;
signal \N__4515\ : std_logic;
signal \N__4502\ : std_logic;
signal \N__4501\ : std_logic;
signal \N__4498\ : std_logic;
signal \N__4497\ : std_logic;
signal \N__4494\ : std_logic;
signal \N__4493\ : std_logic;
signal \N__4492\ : std_logic;
signal \N__4489\ : std_logic;
signal \N__4486\ : std_logic;
signal \N__4485\ : std_logic;
signal \N__4482\ : std_logic;
signal \N__4479\ : std_logic;
signal \N__4476\ : std_logic;
signal \N__4473\ : std_logic;
signal \N__4470\ : std_logic;
signal \N__4467\ : std_logic;
signal \N__4462\ : std_logic;
signal \N__4459\ : std_logic;
signal \N__4458\ : std_logic;
signal \N__4457\ : std_logic;
signal \N__4454\ : std_logic;
signal \N__4447\ : std_logic;
signal \N__4444\ : std_logic;
signal \N__4439\ : std_logic;
signal \N__4430\ : std_logic;
signal \N__4427\ : std_logic;
signal \N__4424\ : std_logic;
signal \N__4421\ : std_logic;
signal \N__4418\ : std_logic;
signal \N__4417\ : std_logic;
signal \N__4414\ : std_logic;
signal \N__4413\ : std_logic;
signal \N__4412\ : std_logic;
signal \N__4411\ : std_logic;
signal \N__4408\ : std_logic;
signal \N__4405\ : std_logic;
signal \N__4402\ : std_logic;
signal \N__4397\ : std_logic;
signal \N__4388\ : std_logic;
signal \N__4387\ : std_logic;
signal \N__4384\ : std_logic;
signal \N__4383\ : std_logic;
signal \N__4380\ : std_logic;
signal \N__4377\ : std_logic;
signal \N__4374\ : std_logic;
signal \N__4369\ : std_logic;
signal \N__4366\ : std_logic;
signal \N__4363\ : std_logic;
signal \N__4358\ : std_logic;
signal \N__4355\ : std_logic;
signal \N__4352\ : std_logic;
signal \N__4351\ : std_logic;
signal \N__4348\ : std_logic;
signal \N__4345\ : std_logic;
signal \N__4340\ : std_logic;
signal \N__4337\ : std_logic;
signal \N__4334\ : std_logic;
signal \N__4331\ : std_logic;
signal \N__4328\ : std_logic;
signal \N__4325\ : std_logic;
signal \N__4322\ : std_logic;
signal \N__4319\ : std_logic;
signal \N__4316\ : std_logic;
signal \N__4313\ : std_logic;
signal \N__4310\ : std_logic;
signal \N__4309\ : std_logic;
signal \N__4308\ : std_logic;
signal \N__4305\ : std_logic;
signal \N__4302\ : std_logic;
signal \N__4299\ : std_logic;
signal \N__4292\ : std_logic;
signal \N__4289\ : std_logic;
signal \N__4286\ : std_logic;
signal \N__4283\ : std_logic;
signal \N__4280\ : std_logic;
signal \N__4277\ : std_logic;
signal \N__4274\ : std_logic;
signal \N__4273\ : std_logic;
signal \N__4272\ : std_logic;
signal \N__4271\ : std_logic;
signal \N__4268\ : std_logic;
signal \N__4267\ : std_logic;
signal \N__4264\ : std_logic;
signal \N__4259\ : std_logic;
signal \N__4256\ : std_logic;
signal \N__4253\ : std_logic;
signal \N__4252\ : std_logic;
signal \N__4251\ : std_logic;
signal \N__4250\ : std_logic;
signal \N__4249\ : std_logic;
signal \N__4248\ : std_logic;
signal \N__4243\ : std_logic;
signal \N__4238\ : std_logic;
signal \N__4233\ : std_logic;
signal \N__4228\ : std_logic;
signal \N__4225\ : std_logic;
signal \N__4214\ : std_logic;
signal \N__4213\ : std_logic;
signal \N__4210\ : std_logic;
signal \N__4207\ : std_logic;
signal \N__4206\ : std_logic;
signal \N__4205\ : std_logic;
signal \N__4204\ : std_logic;
signal \N__4203\ : std_logic;
signal \N__4198\ : std_logic;
signal \N__4195\ : std_logic;
signal \N__4194\ : std_logic;
signal \N__4191\ : std_logic;
signal \N__4188\ : std_logic;
signal \N__4185\ : std_logic;
signal \N__4184\ : std_logic;
signal \N__4183\ : std_logic;
signal \N__4180\ : std_logic;
signal \N__4179\ : std_logic;
signal \N__4176\ : std_logic;
signal \N__4173\ : std_logic;
signal \N__4166\ : std_logic;
signal \N__4161\ : std_logic;
signal \N__4158\ : std_logic;
signal \N__4155\ : std_logic;
signal \N__4150\ : std_logic;
signal \N__4147\ : std_logic;
signal \N__4136\ : std_logic;
signal \N__4135\ : std_logic;
signal \N__4132\ : std_logic;
signal \N__4129\ : std_logic;
signal \N__4126\ : std_logic;
signal \N__4121\ : std_logic;
signal \N__4118\ : std_logic;
signal \N__4117\ : std_logic;
signal \N__4112\ : std_logic;
signal \N__4109\ : std_logic;
signal \N__4106\ : std_logic;
signal \N__4103\ : std_logic;
signal \N__4100\ : std_logic;
signal \N__4097\ : std_logic;
signal \N__4094\ : std_logic;
signal \N__4091\ : std_logic;
signal \N__4088\ : std_logic;
signal \N__4085\ : std_logic;
signal \N__4082\ : std_logic;
signal \N__4079\ : std_logic;
signal \N__4076\ : std_logic;
signal \N__4073\ : std_logic;
signal \N__4070\ : std_logic;
signal \N__4067\ : std_logic;
signal \N__4064\ : std_logic;
signal \N__4061\ : std_logic;
signal \N__4058\ : std_logic;
signal \N__4055\ : std_logic;
signal \N__4052\ : std_logic;
signal \N__4049\ : std_logic;
signal \N__4046\ : std_logic;
signal \N__4043\ : std_logic;
signal \N__4040\ : std_logic;
signal \N__4037\ : std_logic;
signal \N__4034\ : std_logic;
signal \N__4031\ : std_logic;
signal \N__4028\ : std_logic;
signal \N__4025\ : std_logic;
signal \N__4022\ : std_logic;
signal \N__4019\ : std_logic;
signal \N__4016\ : std_logic;
signal \N__4013\ : std_logic;
signal \N__4010\ : std_logic;
signal \N__4009\ : std_logic;
signal \N__4006\ : std_logic;
signal \N__4003\ : std_logic;
signal \N__4000\ : std_logic;
signal \N__3997\ : std_logic;
signal \N__3992\ : std_logic;
signal \N__3989\ : std_logic;
signal \N__3986\ : std_logic;
signal \N__3985\ : std_logic;
signal \N__3982\ : std_logic;
signal \N__3979\ : std_logic;
signal \N__3976\ : std_logic;
signal \N__3971\ : std_logic;
signal \N__3968\ : std_logic;
signal \N__3967\ : std_logic;
signal \N__3966\ : std_logic;
signal \N__3965\ : std_logic;
signal \N__3964\ : std_logic;
signal \N__3963\ : std_logic;
signal \N__3960\ : std_logic;
signal \N__3955\ : std_logic;
signal \N__3952\ : std_logic;
signal \N__3949\ : std_logic;
signal \N__3946\ : std_logic;
signal \N__3943\ : std_logic;
signal \N__3940\ : std_logic;
signal \N__3937\ : std_logic;
signal \N__3926\ : std_logic;
signal \N__3925\ : std_logic;
signal \N__3922\ : std_logic;
signal \N__3919\ : std_logic;
signal \N__3916\ : std_logic;
signal \N__3913\ : std_logic;
signal \N__3912\ : std_logic;
signal \N__3909\ : std_logic;
signal \N__3906\ : std_logic;
signal \N__3903\ : std_logic;
signal \N__3900\ : std_logic;
signal \N__3897\ : std_logic;
signal \N__3890\ : std_logic;
signal \N__3889\ : std_logic;
signal \N__3888\ : std_logic;
signal \N__3885\ : std_logic;
signal \N__3882\ : std_logic;
signal \N__3879\ : std_logic;
signal \N__3876\ : std_logic;
signal \N__3875\ : std_logic;
signal \N__3872\ : std_logic;
signal \N__3869\ : std_logic;
signal \N__3866\ : std_logic;
signal \N__3863\ : std_logic;
signal \N__3860\ : std_logic;
signal \N__3857\ : std_logic;
signal \N__3848\ : std_logic;
signal \N__3845\ : std_logic;
signal \N__3842\ : std_logic;
signal \N__3839\ : std_logic;
signal \N__3836\ : std_logic;
signal \N__3833\ : std_logic;
signal \N__3830\ : std_logic;
signal \N__3827\ : std_logic;
signal \N__3824\ : std_logic;
signal \N__3821\ : std_logic;
signal \N__3820\ : std_logic;
signal \N__3817\ : std_logic;
signal \N__3814\ : std_logic;
signal \N__3809\ : std_logic;
signal \N__3806\ : std_logic;
signal \N__3803\ : std_logic;
signal \N__3800\ : std_logic;
signal \N__3797\ : std_logic;
signal \N__3794\ : std_logic;
signal \N__3791\ : std_logic;
signal \N__3788\ : std_logic;
signal \N__3785\ : std_logic;
signal \N__3782\ : std_logic;
signal \N__3779\ : std_logic;
signal \N__3776\ : std_logic;
signal \N__3773\ : std_logic;
signal \N__3770\ : std_logic;
signal \N__3769\ : std_logic;
signal \N__3766\ : std_logic;
signal \N__3763\ : std_logic;
signal \N__3760\ : std_logic;
signal \N__3757\ : std_logic;
signal \N__3752\ : std_logic;
signal \N__3749\ : std_logic;
signal \N__3746\ : std_logic;
signal \N__3743\ : std_logic;
signal \N__3740\ : std_logic;
signal \N__3737\ : std_logic;
signal \N__3734\ : std_logic;
signal \N__3731\ : std_logic;
signal \N__3728\ : std_logic;
signal \N__3725\ : std_logic;
signal \N__3722\ : std_logic;
signal \N__3719\ : std_logic;
signal \N__3718\ : std_logic;
signal \N__3715\ : std_logic;
signal \N__3712\ : std_logic;
signal \N__3711\ : std_logic;
signal \N__3708\ : std_logic;
signal \N__3705\ : std_logic;
signal \N__3704\ : std_logic;
signal \N__3701\ : std_logic;
signal \N__3700\ : std_logic;
signal \N__3695\ : std_logic;
signal \N__3692\ : std_logic;
signal \N__3689\ : std_logic;
signal \N__3686\ : std_logic;
signal \N__3681\ : std_logic;
signal \N__3678\ : std_logic;
signal \N__3671\ : std_logic;
signal \N__3670\ : std_logic;
signal \N__3667\ : std_logic;
signal \N__3666\ : std_logic;
signal \N__3663\ : std_logic;
signal \N__3662\ : std_logic;
signal \N__3659\ : std_logic;
signal \N__3656\ : std_logic;
signal \N__3653\ : std_logic;
signal \N__3650\ : std_logic;
signal \N__3645\ : std_logic;
signal \N__3644\ : std_logic;
signal \N__3643\ : std_logic;
signal \N__3636\ : std_logic;
signal \N__3631\ : std_logic;
signal \N__3626\ : std_logic;
signal \N__3623\ : std_logic;
signal \N__3622\ : std_logic;
signal \N__3619\ : std_logic;
signal \N__3616\ : std_logic;
signal \N__3611\ : std_logic;
signal \N__3608\ : std_logic;
signal \N__3605\ : std_logic;
signal \N__3602\ : std_logic;
signal \N__3599\ : std_logic;
signal \N__3598\ : std_logic;
signal \N__3593\ : std_logic;
signal \N__3590\ : std_logic;
signal \N__3587\ : std_logic;
signal \N__3584\ : std_logic;
signal \N__3581\ : std_logic;
signal \N__3578\ : std_logic;
signal \N__3575\ : std_logic;
signal \N__3572\ : std_logic;
signal \N__3569\ : std_logic;
signal \N__3566\ : std_logic;
signal \N__3563\ : std_logic;
signal \N__3560\ : std_logic;
signal \N__3557\ : std_logic;
signal \N__3554\ : std_logic;
signal \N__3551\ : std_logic;
signal \N__3548\ : std_logic;
signal \N__3547\ : std_logic;
signal \N__3546\ : std_logic;
signal \N__3545\ : std_logic;
signal \N__3542\ : std_logic;
signal \N__3541\ : std_logic;
signal \N__3538\ : std_logic;
signal \N__3537\ : std_logic;
signal \N__3534\ : std_logic;
signal \N__3527\ : std_logic;
signal \N__3524\ : std_logic;
signal \N__3523\ : std_logic;
signal \N__3520\ : std_logic;
signal \N__3517\ : std_logic;
signal \N__3516\ : std_logic;
signal \N__3515\ : std_logic;
signal \N__3514\ : std_logic;
signal \N__3511\ : std_logic;
signal \N__3508\ : std_logic;
signal \N__3503\ : std_logic;
signal \N__3500\ : std_logic;
signal \N__3493\ : std_logic;
signal \N__3486\ : std_logic;
signal \N__3479\ : std_logic;
signal \N__3476\ : std_logic;
signal \N__3473\ : std_logic;
signal \N__3470\ : std_logic;
signal \N__3467\ : std_logic;
signal \N__3464\ : std_logic;
signal \N__3461\ : std_logic;
signal \N__3458\ : std_logic;
signal \N__3455\ : std_logic;
signal \N__3452\ : std_logic;
signal \N__3449\ : std_logic;
signal \N__3446\ : std_logic;
signal \N__3443\ : std_logic;
signal \N__3440\ : std_logic;
signal \N__3437\ : std_logic;
signal \N__3434\ : std_logic;
signal \N__3433\ : std_logic;
signal \N__3432\ : std_logic;
signal \N__3429\ : std_logic;
signal \N__3428\ : std_logic;
signal \N__3425\ : std_logic;
signal \N__3424\ : std_logic;
signal \N__3421\ : std_logic;
signal \N__3418\ : std_logic;
signal \N__3413\ : std_logic;
signal \N__3410\ : std_logic;
signal \N__3409\ : std_logic;
signal \N__3406\ : std_logic;
signal \N__3401\ : std_logic;
signal \N__3398\ : std_logic;
signal \N__3395\ : std_logic;
signal \N__3386\ : std_logic;
signal \N__3383\ : std_logic;
signal \N__3380\ : std_logic;
signal \N__3377\ : std_logic;
signal \N__3376\ : std_logic;
signal \N__3375\ : std_logic;
signal \N__3374\ : std_logic;
signal \N__3371\ : std_logic;
signal \N__3366\ : std_logic;
signal \N__3363\ : std_logic;
signal \N__3356\ : std_logic;
signal \N__3355\ : std_logic;
signal \N__3352\ : std_logic;
signal \N__3351\ : std_logic;
signal \N__3348\ : std_logic;
signal \N__3345\ : std_logic;
signal \N__3340\ : std_logic;
signal \N__3335\ : std_logic;
signal \N__3332\ : std_logic;
signal \N__3329\ : std_logic;
signal \N__3328\ : std_logic;
signal \N__3327\ : std_logic;
signal \N__3324\ : std_logic;
signal \N__3319\ : std_logic;
signal \N__3314\ : std_logic;
signal \N__3311\ : std_logic;
signal \N__3308\ : std_logic;
signal \N__3305\ : std_logic;
signal \N__3302\ : std_logic;
signal \N__3301\ : std_logic;
signal \N__3298\ : std_logic;
signal \N__3297\ : std_logic;
signal \N__3296\ : std_logic;
signal \N__3295\ : std_logic;
signal \N__3292\ : std_logic;
signal \N__3289\ : std_logic;
signal \N__3286\ : std_logic;
signal \N__3281\ : std_logic;
signal \N__3272\ : std_logic;
signal \N__3269\ : std_logic;
signal \N__3268\ : std_logic;
signal \N__3267\ : std_logic;
signal \N__3266\ : std_logic;
signal \N__3265\ : std_logic;
signal \N__3262\ : std_logic;
signal \N__3255\ : std_logic;
signal \N__3252\ : std_logic;
signal \N__3245\ : std_logic;
signal \N__3242\ : std_logic;
signal \N__3239\ : std_logic;
signal \N__3236\ : std_logic;
signal \N__3233\ : std_logic;
signal \N__3230\ : std_logic;
signal \N__3227\ : std_logic;
signal \N__3224\ : std_logic;
signal \N__3221\ : std_logic;
signal \N__3218\ : std_logic;
signal \N__3215\ : std_logic;
signal \N__3212\ : std_logic;
signal \N__3211\ : std_logic;
signal \N__3210\ : std_logic;
signal \N__3207\ : std_logic;
signal \N__3202\ : std_logic;
signal \N__3197\ : std_logic;
signal \N__3194\ : std_logic;
signal \N__3191\ : std_logic;
signal \N__3188\ : std_logic;
signal \N__3185\ : std_logic;
signal \N__3184\ : std_logic;
signal \N__3183\ : std_logic;
signal \N__3182\ : std_logic;
signal \N__3181\ : std_logic;
signal \N__3180\ : std_logic;
signal \N__3177\ : std_logic;
signal \N__3172\ : std_logic;
signal \N__3167\ : std_logic;
signal \N__3164\ : std_logic;
signal \N__3155\ : std_logic;
signal \N__3154\ : std_logic;
signal \N__3153\ : std_logic;
signal \N__3152\ : std_logic;
signal \N__3151\ : std_logic;
signal \N__3148\ : std_logic;
signal \N__3145\ : std_logic;
signal \N__3140\ : std_logic;
signal \N__3137\ : std_logic;
signal \N__3132\ : std_logic;
signal \N__3127\ : std_logic;
signal \N__3124\ : std_logic;
signal \N__3119\ : std_logic;
signal \N__3116\ : std_logic;
signal \N__3113\ : std_logic;
signal \N__3110\ : std_logic;
signal \N__3107\ : std_logic;
signal \N__3106\ : std_logic;
signal \N__3103\ : std_logic;
signal \N__3100\ : std_logic;
signal \N__3097\ : std_logic;
signal \N__3092\ : std_logic;
signal \N__3089\ : std_logic;
signal \N__3086\ : std_logic;
signal \N__3083\ : std_logic;
signal \N__3080\ : std_logic;
signal \N__3077\ : std_logic;
signal \N__3074\ : std_logic;
signal \N__3071\ : std_logic;
signal \N__3068\ : std_logic;
signal \N__3065\ : std_logic;
signal \N__3062\ : std_logic;
signal \N__3059\ : std_logic;
signal \N__3056\ : std_logic;
signal \N__3053\ : std_logic;
signal \N__3050\ : std_logic;
signal \N__3047\ : std_logic;
signal \N__3044\ : std_logic;
signal \N__3041\ : std_logic;
signal \N__3038\ : std_logic;
signal \N__3035\ : std_logic;
signal \N__3032\ : std_logic;
signal \N__3029\ : std_logic;
signal \N__3026\ : std_logic;
signal \N__3023\ : std_logic;
signal \N__3020\ : std_logic;
signal \N__3017\ : std_logic;
signal \N__3014\ : std_logic;
signal \N__3011\ : std_logic;
signal \N__3008\ : std_logic;
signal \N__3007\ : std_logic;
signal \N__3002\ : std_logic;
signal \N__2999\ : std_logic;
signal \N__2998\ : std_logic;
signal \N__2995\ : std_logic;
signal \N__2992\ : std_logic;
signal \N__2989\ : std_logic;
signal \N__2984\ : std_logic;
signal \N__2981\ : std_logic;
signal \N__2978\ : std_logic;
signal \N__2975\ : std_logic;
signal \N__2972\ : std_logic;
signal \N__2969\ : std_logic;
signal \N__2966\ : std_logic;
signal \N__2963\ : std_logic;
signal \N__2960\ : std_logic;
signal \N__2957\ : std_logic;
signal \N__2954\ : std_logic;
signal \N__2951\ : std_logic;
signal \N__2948\ : std_logic;
signal \N__2945\ : std_logic;
signal \N__2942\ : std_logic;
signal \N__2939\ : std_logic;
signal \N__2936\ : std_logic;
signal \N__2933\ : std_logic;
signal \N__2930\ : std_logic;
signal \N__2927\ : std_logic;
signal \N__2924\ : std_logic;
signal \N__2921\ : std_logic;
signal \N__2918\ : std_logic;
signal \N__2915\ : std_logic;
signal \N__2912\ : std_logic;
signal \N__2909\ : std_logic;
signal \N__2906\ : std_logic;
signal \N__2903\ : std_logic;
signal \N__2900\ : std_logic;
signal \N__2897\ : std_logic;
signal \N__2894\ : std_logic;
signal \N__2891\ : std_logic;
signal \N__2888\ : std_logic;
signal \N__2885\ : std_logic;
signal \N__2882\ : std_logic;
signal \N__2879\ : std_logic;
signal \N__2876\ : std_logic;
signal \N__2873\ : std_logic;
signal \N__2870\ : std_logic;
signal \N__2867\ : std_logic;
signal \N__2864\ : std_logic;
signal \N__2861\ : std_logic;
signal \N__2858\ : std_logic;
signal \N__2855\ : std_logic;
signal \N__2852\ : std_logic;
signal \N__2849\ : std_logic;
signal \GNDG0\ : std_logic;
signal \VCCG0\ : std_logic;
signal \INVseq.counter.T_0_2_rep1C_net\ : std_logic;
signal clk_c : std_logic;
signal buf_clk_1 : std_logic;
signal \pc.N_21_0_cascade_\ : std_logic;
signal \seq_D_6_cascade_\ : std_logic;
signal \pc.G_12_i_a3_1\ : std_logic;
signal \pc.program_counter_m_3_cascade_\ : std_logic;
signal \pc.tbuf.gZ0Z3\ : std_logic;
signal \pc.tbuf.g0Z0Z_3_cascade_\ : std_logic;
signal \bus_3_cascade_\ : std_logic;
signal \INVAR.ff4.qC_net\ : std_logic;
signal \seq_MAR_LD_1_0\ : std_logic;
signal \pc.program_counter_m_3\ : std_logic;
signal \seq.DZ0Z_0_cascade_\ : std_logic;
signal \seq_un1_IR_OE_4_1_cascade_\ : std_logic;
signal \pc.program_counter_RNO_5Z0Z_0\ : std_logic;
signal \seq.un17_IR_OE_cascade_\ : std_logic;
signal \seq_PC_LD_0_0_cascade_\ : std_logic;
signal \seq.D_6_x\ : std_logic;
signal \INVIR.ff5.q_0_rep1C_net\ : std_logic;
signal \bus_6_cascade_\ : std_logic;
signal \N_5_0_cascade_\ : std_logic;
signal \INVIR.ff7.q_ret_1C_net\ : std_logic;
signal \INVIR.ff5.q_0_nerC_net\ : std_logic;
signal \INVseq.counter.T_4C_net\ : std_logic;
signal \mem_data_2_7_0__g1\ : std_logic;
signal \pc.program_counter_m_0_2_cascade_\ : std_logic;
signal \AR_out_2\ : std_logic;
signal \INVAR.ff3.qC_net\ : std_logic;
signal \AR_out_0\ : std_logic;
signal \mem_data_2_7_0__N_7_0\ : std_logic;
signal \pc.program_counter_m_0_0\ : std_logic;
signal \pc.out_1_2_iv_0_cascade_\ : std_logic;
signal \pc.tbuf.g0Z0Z_1_cascade_\ : std_logic;
signal bus_0 : std_logic;
signal \mem_data_2_7_0__N_14_0\ : std_logic;
signal \ALU_main.N_48_cascade_\ : std_logic;
signal \alu_out_m_7_cascade_\ : std_logic;
signal \acc_out_m_7_cascade_\ : std_logic;
signal out_c_7 : std_logic;
signal \INVout_reg.ff8.qC_net\ : std_logic;
signal \pc.out_1_2_iv_0\ : std_logic;
signal \pc.program_counter_RNO_7Z0Z_0_cascade_\ : std_logic;
signal \pc.program_counter_RNO_3Z0Z_0\ : std_logic;
signal \pc.program_counter_RNO_8Z0Z_0\ : std_logic;
signal \INVmar.ff1.q_nerC_net\ : std_logic;
signal \ROM_OE_cascade_\ : std_logic;
signal \pc.program_counter_m_2\ : std_logic;
signal \pc.out_1_0_iv_0\ : std_logic;
signal \pc.G_10_0_a11_2_1_cascade_\ : std_logic;
signal \pc.N_23\ : std_logic;
signal \pc.program_counter_RNO_6Z0Z_2_cascade_\ : std_logic;
signal \pc.G_10_0_a11_5_2\ : std_logic;
signal \seq.S1_1Z0Z_0_cascade_\ : std_logic;
signal \seq_S1_0_cascade_\ : std_logic;
signal \pc.N_16\ : std_logic;
signal bus_6 : std_logic;
signal ir_out_fast_4 : std_logic;
signal \seq.counter.T_RNI0T6TZ0Z_4_cascade_\ : std_logic;
signal ir_out_7_rep1 : std_logic;
signal \INVIR.ff7.q_0_fastC_net\ : std_logic;
signal \seq_T_2_rep1\ : std_logic;
signal \seq.D_1_0_x_cascade_\ : std_logic;
signal \INVIR.ff6.q_ret_1C_net\ : std_logic;
signal \seq.B_LD_0_2_tz_cascade_\ : std_logic;
signal \seq.counter.T_RNIR83I4_0Z0Z_3\ : std_logic;
signal \IR_ff6_q_0_fast\ : std_logic;
signal \IR_ff7_q_ret_1_fast\ : std_logic;
signal \seq.counter.T_0_fast_RNIP4D21Z0Z_2_cascade_\ : std_logic;
signal \T_0_fast_RNILB791_2_cascade_\ : std_logic;
signal \pc.G_12_i_0\ : std_logic;
signal \seq.counter.T_0_fast_RNIG89VZ0Z_2_cascade_\ : std_logic;
signal ir_out_fast_7 : std_logic;
signal \INVseq.counter.T_0_fast_2C_net\ : std_logic;
signal \seq.S0_0_i_N_3LZ0Z3\ : std_logic;
signal ir_out_i_2_6 : std_logic;
signal \INVIR.ff7.q_0_nerC_net\ : std_logic;
signal \seq.counter.T_fast_2\ : std_logic;
signal \seq_un1_IR_OE_4_1\ : std_logic;
signal \g0_0_1_cascade_\ : std_logic;
signal \seq.counter.un7_ACC_LD_0\ : std_logic;
signal \seq.un1_ALU_en_0Z0Z_1\ : std_logic;
signal \seq.counter.un7_ACC_LD_0_cascade_\ : std_logic;
signal \IR_OE_2_cascade_\ : std_logic;
signal bus_2 : std_logic;
signal \seq.g2Z0Z_0\ : std_logic;
signal \IR_OE_1_cascade_\ : std_logic;
signal \pc.un1_inc_0\ : std_logic;
signal \pc.G_12_i_a3_2_3\ : std_logic;
signal \pc.G_12_i_a3_2_1\ : std_logic;
signal \seq.counter.T8_1_cascade_\ : std_logic;
signal \pc.g1_0\ : std_logic;
signal \pc.N_188_0\ : std_logic;
signal \seq_T_0\ : std_logic;
signal \INVseq.counter.T_0C_net\ : std_logic;
signal \N_30\ : std_logic;
signal \pc.G_10_0_1_0_cascade_\ : std_logic;
signal \pc.G_10_0_sx\ : std_logic;
signal \pc.G_10_0_5_1\ : std_logic;
signal \ALU_main_N_43_0\ : std_logic;
signal \pc.program_counterZ0Z_2\ : std_logic;
signal \pc.program_counterZ0Z_0\ : std_logic;
signal \seq_S0_0_i\ : std_logic;
signal \bfn_4_12_0_\ : std_logic;
signal \ALU_main.un1_A_cry_0_c_THRU_CO\ : std_logic;
signal \ALU_main.un1_A_cry_0\ : std_logic;
signal \ALU_main.un1_A_axb_2_l_ofxZ0\ : std_logic;
signal \un1_A_cry_1_c_RNITKPO2\ : std_logic;
signal \ALU_main.un1_A_cry_1\ : std_logic;
signal \ALU_main.un1_A_cry_2\ : std_logic;
signal \ALU_main.un1_A_cry_3\ : std_logic;
signal \ALU_main.un1_A_cry_4\ : std_logic;
signal \ALU_main.un1_A_cry_5\ : std_logic;
signal \ALU_main.un1_A_cry_6\ : std_logic;
signal \bfn_4_13_0_\ : std_logic;
signal \ALU_main.un1_A_cry_6_c_RNIP89EZ0Z2\ : std_logic;
signal \ALU_main.un1_A_cry_5_c_RNIDLAPZ0Z2\ : std_logic;
signal \ALU_main_N_44_0_cascade_\ : std_logic;
signal \un1_A_cry_2_c_RNI1TTO2\ : std_logic;
signal \pc.N_10_i\ : std_logic;
signal \pc.G_10_0_1_1\ : std_logic;
signal \pc.G_10_0_1\ : std_logic;
signal \ALU_main_N_44_1\ : std_logic;
signal \pc.un1_inc_0_0\ : std_logic;
signal \pc.out_1_iv_1_1\ : std_logic;
signal \mem_data_2_7_0__N_16_0\ : std_logic;
signal \pc.g0_rn_1\ : std_logic;
signal \pc.g0_sn_cascade_\ : std_logic;
signal alu_out_m_0_3 : std_logic;
signal \pc.program_counterZ0Z_3\ : std_logic;
signal \seq_un1_AR_OE_0_0\ : std_logic;
signal ir_out_6 : std_logic;
signal \AR.ff4.AR_out_3\ : std_logic;
signal ir_out_3 : std_logic;
signal \pc.tbuf.g0_0_1_0\ : std_logic;
signal \AR_out_m_3_cascade_\ : std_logic;
signal \pc.g0_0\ : std_logic;
signal ir_out_5 : std_logic;
signal bus_7 : std_logic;
signal \N_5_0\ : std_logic;
signal \N_1_0_cascade_\ : std_logic;
signal \seq_un1_HLT_0\ : std_logic;
signal \INVseq.q_ret_1C_net\ : std_logic;
signal \seq.un1_HLT_1_reti\ : std_logic;
signal \N_2_0\ : std_logic;
signal \seq.un1_HLT_1\ : std_logic;
signal \INVseq.q_retC_net\ : std_logic;
signal \bus_1_cascade_\ : std_logic;
signal \seq_D_6\ : std_logic;
signal \T_0_fast_RNILB791_2\ : std_logic;
signal \AR_out_1\ : std_logic;
signal \INVAR.ff2.qC_net\ : std_logic;
signal \seq.D_3\ : std_logic;
signal \seq.counter.ACC_LD_0_0_cascade_\ : std_logic;
signal \pc.program_counter_m_0_1\ : std_logic;
signal \pc.tbuf.out_1_1_ivZ0Z_0\ : std_logic;
signal \mem_data_2_7_0__N_11_0_cascade_\ : std_logic;
signal \pc.program_counter_4_rn_2_1\ : std_logic;
signal \pc.program_counter_4_sn_1\ : std_logic;
signal \pc.g0_1_0_cascade_\ : std_logic;
signal \pc.program_counterZ0Z_1\ : std_logic;
signal buf_clk_1_g : std_logic;
signal \seq_T_2\ : std_logic;
signal \seq_PC_LD_0_0\ : std_logic;
signal \seq_MAR_LD_2\ : std_logic;
signal \seq.gZ0Z2\ : std_logic;
signal \ALU_main_N_42_0_cascade_\ : std_logic;
signal \un1_A_cry_0_c_RNIPCLO2\ : std_logic;
signal \ALU_main_N_41_0_cascade_\ : std_logic;
signal \un1_A_cry_0_s\ : std_logic;
signal \seq.D_4\ : std_logic;
signal \seq.DZ0Z_0\ : std_logic;
signal \seq.g2Z0Z_1\ : std_logic;
signal \ALU_main.un1_A_axb_0_l_ofxZ0\ : std_logic;
signal \ALU_main.un1_A_axb_3_l_ofxZ0\ : std_logic;
signal \ALU_main.un1_A_cry_4_c_RNI9D6PZ0Z2\ : std_logic;
signal \ALU_main.N_46_cascade_\ : std_logic;
signal ir_out_i_2_5 : std_logic;
signal ir_out_4_rep1 : std_logic;
signal \IR_ff7_q_0_fast\ : std_logic;
signal \seq.counter.TZ0Z_4\ : std_logic;
signal ir_out_7 : std_logic;
signal \seq.g0_i_a3_0Z0Z_2_cascade_\ : std_logic;
signal \seq.g0_i_a3Z0Z_2\ : std_logic;
signal \seq_S0_0_cascade_\ : std_logic;
signal \ALU_main.un1_A_axb_5_l_ofxZ0\ : std_logic;
signal \seq.counter.TZ0Z_3\ : std_logic;
signal \seq.D_2\ : std_logic;
signal \seq.B_LD_0_2_tz\ : std_logic;
signal \seq.D_1\ : std_logic;
signal \ALU_main.un1_A_axb_1_l_ofxZ0\ : std_logic;
signal \INVb_reg.ff5.qC_net\ : std_logic;
signal \ALU_main.un1_A_axb_4_l_ofxZ0\ : std_logic;
signal \ALU_main.N_47\ : std_logic;
signal acc_out_6 : std_logic;
signal \ALU_main.un1_A_axb_6_l_ofxZ0\ : std_logic;
signal acc_out_7 : std_logic;
signal acc_out_5 : std_logic;
signal acc_out_3 : std_logic;
signal \INVacc.ff7.qC_net\ : std_logic;
signal \ALU_main.un1_A_cry_3_c_RNI552PZ0Z2\ : std_logic;
signal \seq_un1_ALU_en_0\ : std_logic;
signal \seq_S1_0\ : std_logic;
signal \alu_out_m_4_cascade_\ : std_logic;
signal bus_4 : std_logic;
signal \bus_4_cascade_\ : std_logic;
signal ir_out_4 : std_logic;
signal \N_4_0\ : std_logic;
signal b_reg_out_4 : std_logic;
signal \seq_S0_0\ : std_logic;
signal \ALU_main.N_45\ : std_logic;
signal bus_5 : std_logic;
signal \INVIR.ff2.q_nerC_net\ : std_logic;
signal acc_out_0 : std_logic;
signal acc_out_1 : std_logic;
signal acc_out_2 : std_logic;
signal \INVacc.ff1.qC_net\ : std_logic;
signal \seq_ACC_LD_0_i\ : std_logic;
signal \INVmar.ff4.q_nerC_net\ : std_logic;
signal \mar.MAR_LD_0_0\ : std_logic;
signal b_reg_out_5 : std_logic;
signal acc_out_m_7 : std_logic;
signal alu_out_m_7 : std_logic;
signal b_reg_out_7 : std_logic;
signal b_reg_out_0 : std_logic;
signal \INVb_reg.ff6.qC_net\ : std_logic;
signal \mem.i2_mux_cascade_\ : std_logic;
signal \pc.N_7\ : std_logic;
signal \mem_data_2_7_0__N_29_mux_cascade_\ : std_logic;
signal out_c_6 : std_logic;
signal \INVout_reg.ff7.qC_net\ : std_logic;
signal mar_out_2 : std_logic;
signal mar_out_1 : std_logic;
signal mar_out_3 : std_logic;
signal mar_out_0 : std_logic;
signal \mem_data_2_7_0__i2_mux_0\ : std_logic;
signal b_reg_out_1 : std_logic;
signal acc_out_m_6 : std_logic;
signal alu_out_m_6 : std_logic;
signal \mem_data_2_7_0__N_29_mux\ : std_logic;
signal b_reg_out_6 : std_logic;
signal \INVb_reg.ff2.qC_net\ : std_logic;
signal acc_out_m_5 : std_logic;
signal alu_out_m_5 : std_logic;
signal m20 : std_logic;
signal \ROM_OE\ : std_logic;
signal out_c_5 : std_logic;
signal \INVout_reg.ff6.qC_net\ : std_logic;
signal out_c_2 : std_logic;
signal out_c_0 : std_logic;
signal \INVout_reg.ff3.qC_net\ : std_logic;
signal \pc.tbuf.g0Z0Z_1\ : std_logic;
signal \IR_OE_0\ : std_logic;
signal alu_out_m_0_0 : std_logic;
signal ir_out_0 : std_logic;
signal \INVIR.ff1.q_nerC_net\ : std_logic;
signal inc : std_logic;
signal alu_out_m_0_2 : std_logic;
signal ir_out_2 : std_logic;
signal \IR_OE_2\ : std_logic;
signal \pc.tbuf.g0_1_1\ : std_logic;
signal b_reg_out_2 : std_logic;
signal \INVb_reg.ff3.qC_net\ : std_logic;
signal \IR_OE_1\ : std_logic;
signal \pc.g0_1_0\ : std_logic;
signal ir_out_1 : std_logic;
signal alu_out_m_0_1 : std_logic;
signal out_c_1 : std_logic;
signal alu_out_m_4 : std_logic;
signal \mem_data_2_7_0__i2_mux_i_m\ : std_logic;
signal acc_out_4 : std_logic;
signal out_c_4 : std_logic;
signal \INVout_reg.ff2.qC_net\ : std_logic;
signal b_reg_out_3 : std_logic;
signal \INVb_reg.ff4.qC_net\ : std_logic;
signal \seq_B_LD_0_i\ : std_logic;
signal \pc.tbuf.g0_0_0\ : std_logic;
signal \pc.tbuf.g0Z0Z_3\ : std_logic;
signal \pc.tbuf.gZ0Z2\ : std_logic;
signal alu_out_m_1_3 : std_logic;
signal out_c_3 : std_logic;
signal \_gnd_net_\ : std_logic;
signal \INVout_reg.ff4.qC_net\ : std_logic;
signal \OUT_LD\ : std_logic;
signal clr_c_g : std_logic;

signal clr_wire : std_logic;
signal out_wire : std_logic_vector(7 downto 0);
signal clk_wire : std_logic;

begin
    clr_wire <= clr;
    out <= out_wire;
    clk_wire <= clk;

    \clr_ibuf_gb_io_preiogbuf\ : PRE_IO_GBUF
    port map (
            PADSIGNALTOGLOBALBUFFER => \N__9027\,
            GLOBALBUFFEROUTPUT => clr_c_g
        );

    \clr_ibuf_gb_io_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9029\,
            DIN => \N__9028\,
            DOUT => \N__9027\,
            PACKAGEPIN => clr_wire
        );

    \clr_ibuf_gb_io_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__9029\,
            PADOUT => \N__9028\,
            PADIN => \N__9027\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \out_obuf_7_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__9018\,
            DIN => \N__9017\,
            DOUT => \N__9016\,
            PACKAGEPIN => out_wire(7)
        );

    \out_obuf_7_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9018\,
            PADOUT => \N__9017\,
            PADIN => \N__9016\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__3047\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \out_obuf_4_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9009\,
            DIN => \N__9008\,
            DOUT => \N__9007\,
            PACKAGEPIN => out_wire(4)
        );

    \out_obuf_4_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9009\,
            PADOUT => \N__9008\,
            PADIN => \N__9007\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7844\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \out_obuf_3_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__9000\,
            DIN => \N__8999\,
            DOUT => \N__8998\,
            PACKAGEPIN => out_wire(3)
        );

    \out_obuf_3_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__9000\,
            PADOUT => \N__8999\,
            PADIN => \N__8998\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7493\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \out_obuf_6_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8991\,
            DIN => \N__8990\,
            DOUT => \N__8989\,
            PACKAGEPIN => out_wire(6)
        );

    \out_obuf_6_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8991\,
            PADOUT => \N__8990\,
            PADIN => \N__8989\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__7205\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \out_obuf_5_iopad\ : IO_PAD
    generic map (
            IO_STANDARD => "SB_LVCMOS",
            PULLUP => '0'
        )
    port map (
            OE => \N__8982\,
            DIN => \N__8981\,
            DOUT => \N__8980\,
            PACKAGEPIN => out_wire(5)
        );

    \out_obuf_5_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8982\,
            PADOUT => \N__8981\,
            PADIN => \N__8980\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6422\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \out_obuf_0_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8973\,
            DIN => \N__8972\,
            DOUT => \N__8971\,
            PACKAGEPIN => out_wire(0)
        );

    \out_obuf_0_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8973\,
            PADOUT => \N__8972\,
            PADIN => \N__8971\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6398\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \clk_ibuf_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8964\,
            DIN => \N__8963\,
            DOUT => \N__8962\,
            PACKAGEPIN => clk_wire
        );

    \clk_ibuf_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "000001"
        )
    port map (
            PADOEN => \N__8964\,
            PADOUT => \N__8963\,
            PADIN => \N__8962\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => clk_c,
            DOUT0 => '0',
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \out_obuf_2_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8955\,
            DIN => \N__8954\,
            DOUT => \N__8953\,
            PACKAGEPIN => out_wire(2)
        );

    \out_obuf_2_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8955\,
            PADOUT => \N__8954\,
            PADIN => \N__8953\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__6407\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \out_obuf_1_iopad\ : IO_PAD
    generic map (
            PULLUP => '0',
            IO_STANDARD => "SB_LVCMOS"
        )
    port map (
            OE => \N__8946\,
            DIN => \N__8945\,
            DOUT => \N__8944\,
            PACKAGEPIN => out_wire(1)
        );

    \out_obuf_1_preio\ : PRE_IO
    generic map (
            NEG_TRIGGER => '0',
            PIN_TYPE => "011001"
        )
    port map (
            PADOEN => \N__8946\,
            PADOUT => \N__8945\,
            PADIN => \N__8944\,
            CLOCKENABLE => 'H',
            DOUT1 => '0',
            OUTPUTENABLE => '0',
            DIN0 => OPEN,
            DOUT0 => \N__8012\,
            INPUTCLK => '0',
            LATCHINPUTVALUE => '0',
            DIN1 => OPEN,
            OUTPUTCLK => '0'
        );

    \I__2290\ : InMux
    port map (
            O => \N__8927\,
            I => \N__8923\
        );

    \I__2289\ : InMux
    port map (
            O => \N__8926\,
            I => \N__8920\
        );

    \I__2288\ : LocalMux
    port map (
            O => \N__8923\,
            I => \N__8916\
        );

    \I__2287\ : LocalMux
    port map (
            O => \N__8920\,
            I => \N__8913\
        );

    \I__2286\ : InMux
    port map (
            O => \N__8919\,
            I => \N__8910\
        );

    \I__2285\ : Span4Mux_v
    port map (
            O => \N__8916\,
            I => \N__8901\
        );

    \I__2284\ : Span4Mux_h
    port map (
            O => \N__8913\,
            I => \N__8901\
        );

    \I__2283\ : LocalMux
    port map (
            O => \N__8910\,
            I => \N__8901\
        );

    \I__2282\ : InMux
    port map (
            O => \N__8909\,
            I => \N__8898\
        );

    \I__2281\ : InMux
    port map (
            O => \N__8908\,
            I => \N__8895\
        );

    \I__2280\ : Span4Mux_h
    port map (
            O => \N__8901\,
            I => \N__8892\
        );

    \I__2279\ : LocalMux
    port map (
            O => \N__8898\,
            I => \N__8889\
        );

    \I__2278\ : LocalMux
    port map (
            O => \N__8895\,
            I => \N__8886\
        );

    \I__2277\ : Odrv4
    port map (
            O => \N__8892\,
            I => \pc.tbuf.g0Z0Z_1\
        );

    \I__2276\ : Odrv12
    port map (
            O => \N__8889\,
            I => \pc.tbuf.g0Z0Z_1\
        );

    \I__2275\ : Odrv4
    port map (
            O => \N__8886\,
            I => \pc.tbuf.g0Z0Z_1\
        );

    \I__2274\ : CascadeMux
    port map (
            O => \N__8879\,
            I => \N__8874\
        );

    \I__2273\ : CascadeMux
    port map (
            O => \N__8878\,
            I => \N__8870\
        );

    \I__2272\ : InMux
    port map (
            O => \N__8877\,
            I => \N__8867\
        );

    \I__2271\ : InMux
    port map (
            O => \N__8874\,
            I => \N__8864\
        );

    \I__2270\ : InMux
    port map (
            O => \N__8873\,
            I => \N__8861\
        );

    \I__2269\ : InMux
    port map (
            O => \N__8870\,
            I => \N__8857\
        );

    \I__2268\ : LocalMux
    port map (
            O => \N__8867\,
            I => \N__8854\
        );

    \I__2267\ : LocalMux
    port map (
            O => \N__8864\,
            I => \N__8849\
        );

    \I__2266\ : LocalMux
    port map (
            O => \N__8861\,
            I => \N__8849\
        );

    \I__2265\ : CascadeMux
    port map (
            O => \N__8860\,
            I => \N__8845\
        );

    \I__2264\ : LocalMux
    port map (
            O => \N__8857\,
            I => \N__8842\
        );

    \I__2263\ : Span4Mux_v
    port map (
            O => \N__8854\,
            I => \N__8839\
        );

    \I__2262\ : Span4Mux_v
    port map (
            O => \N__8849\,
            I => \N__8836\
        );

    \I__2261\ : InMux
    port map (
            O => \N__8848\,
            I => \N__8833\
        );

    \I__2260\ : InMux
    port map (
            O => \N__8845\,
            I => \N__8830\
        );

    \I__2259\ : Span4Mux_s2_h
    port map (
            O => \N__8842\,
            I => \N__8825\
        );

    \I__2258\ : Span4Mux_s2_h
    port map (
            O => \N__8839\,
            I => \N__8825\
        );

    \I__2257\ : Odrv4
    port map (
            O => \N__8836\,
            I => \IR_OE_0\
        );

    \I__2256\ : LocalMux
    port map (
            O => \N__8833\,
            I => \IR_OE_0\
        );

    \I__2255\ : LocalMux
    port map (
            O => \N__8830\,
            I => \IR_OE_0\
        );

    \I__2254\ : Odrv4
    port map (
            O => \N__8825\,
            I => \IR_OE_0\
        );

    \I__2253\ : InMux
    port map (
            O => \N__8816\,
            I => \N__8811\
        );

    \I__2252\ : InMux
    port map (
            O => \N__8815\,
            I => \N__8808\
        );

    \I__2251\ : InMux
    port map (
            O => \N__8814\,
            I => \N__8804\
        );

    \I__2250\ : LocalMux
    port map (
            O => \N__8811\,
            I => \N__8799\
        );

    \I__2249\ : LocalMux
    port map (
            O => \N__8808\,
            I => \N__8799\
        );

    \I__2248\ : InMux
    port map (
            O => \N__8807\,
            I => \N__8796\
        );

    \I__2247\ : LocalMux
    port map (
            O => \N__8804\,
            I => \N__8791\
        );

    \I__2246\ : Span4Mux_v
    port map (
            O => \N__8799\,
            I => \N__8788\
        );

    \I__2245\ : LocalMux
    port map (
            O => \N__8796\,
            I => \N__8785\
        );

    \I__2244\ : InMux
    port map (
            O => \N__8795\,
            I => \N__8782\
        );

    \I__2243\ : InMux
    port map (
            O => \N__8794\,
            I => \N__8779\
        );

    \I__2242\ : Span4Mux_h
    port map (
            O => \N__8791\,
            I => \N__8776\
        );

    \I__2241\ : Odrv4
    port map (
            O => \N__8788\,
            I => alu_out_m_0_0
        );

    \I__2240\ : Odrv4
    port map (
            O => \N__8785\,
            I => alu_out_m_0_0
        );

    \I__2239\ : LocalMux
    port map (
            O => \N__8782\,
            I => alu_out_m_0_0
        );

    \I__2238\ : LocalMux
    port map (
            O => \N__8779\,
            I => alu_out_m_0_0
        );

    \I__2237\ : Odrv4
    port map (
            O => \N__8776\,
            I => alu_out_m_0_0
        );

    \I__2236\ : CascadeMux
    port map (
            O => \N__8765\,
            I => \N__8760\
        );

    \I__2235\ : InMux
    port map (
            O => \N__8764\,
            I => \N__8757\
        );

    \I__2234\ : InMux
    port map (
            O => \N__8763\,
            I => \N__8752\
        );

    \I__2233\ : InMux
    port map (
            O => \N__8760\,
            I => \N__8749\
        );

    \I__2232\ : LocalMux
    port map (
            O => \N__8757\,
            I => \N__8745\
        );

    \I__2231\ : InMux
    port map (
            O => \N__8756\,
            I => \N__8742\
        );

    \I__2230\ : CascadeMux
    port map (
            O => \N__8755\,
            I => \N__8739\
        );

    \I__2229\ : LocalMux
    port map (
            O => \N__8752\,
            I => \N__8736\
        );

    \I__2228\ : LocalMux
    port map (
            O => \N__8749\,
            I => \N__8733\
        );

    \I__2227\ : CascadeMux
    port map (
            O => \N__8748\,
            I => \N__8728\
        );

    \I__2226\ : Span4Mux_v
    port map (
            O => \N__8745\,
            I => \N__8723\
        );

    \I__2225\ : LocalMux
    port map (
            O => \N__8742\,
            I => \N__8723\
        );

    \I__2224\ : InMux
    port map (
            O => \N__8739\,
            I => \N__8720\
        );

    \I__2223\ : Span4Mux_v
    port map (
            O => \N__8736\,
            I => \N__8715\
        );

    \I__2222\ : Span4Mux_s2_h
    port map (
            O => \N__8733\,
            I => \N__8715\
        );

    \I__2221\ : InMux
    port map (
            O => \N__8732\,
            I => \N__8712\
        );

    \I__2220\ : InMux
    port map (
            O => \N__8731\,
            I => \N__8709\
        );

    \I__2219\ : InMux
    port map (
            O => \N__8728\,
            I => \N__8706\
        );

    \I__2218\ : Span4Mux_h
    port map (
            O => \N__8723\,
            I => \N__8703\
        );

    \I__2217\ : LocalMux
    port map (
            O => \N__8720\,
            I => \N__8698\
        );

    \I__2216\ : Span4Mux_h
    port map (
            O => \N__8715\,
            I => \N__8698\
        );

    \I__2215\ : LocalMux
    port map (
            O => \N__8712\,
            I => ir_out_0
        );

    \I__2214\ : LocalMux
    port map (
            O => \N__8709\,
            I => ir_out_0
        );

    \I__2213\ : LocalMux
    port map (
            O => \N__8706\,
            I => ir_out_0
        );

    \I__2212\ : Odrv4
    port map (
            O => \N__8703\,
            I => ir_out_0
        );

    \I__2211\ : Odrv4
    port map (
            O => \N__8698\,
            I => ir_out_0
        );

    \I__2210\ : CEMux
    port map (
            O => \N__8687\,
            I => \N__8680\
        );

    \I__2209\ : CascadeMux
    port map (
            O => \N__8686\,
            I => \N__8669\
        );

    \I__2208\ : CascadeMux
    port map (
            O => \N__8685\,
            I => \N__8656\
        );

    \I__2207\ : CascadeMux
    port map (
            O => \N__8684\,
            I => \N__8651\
        );

    \I__2206\ : CEMux
    port map (
            O => \N__8683\,
            I => \N__8648\
        );

    \I__2205\ : LocalMux
    port map (
            O => \N__8680\,
            I => \N__8645\
        );

    \I__2204\ : CEMux
    port map (
            O => \N__8679\,
            I => \N__8642\
        );

    \I__2203\ : CEMux
    port map (
            O => \N__8678\,
            I => \N__8639\
        );

    \I__2202\ : InMux
    port map (
            O => \N__8677\,
            I => \N__8636\
        );

    \I__2201\ : InMux
    port map (
            O => \N__8676\,
            I => \N__8633\
        );

    \I__2200\ : InMux
    port map (
            O => \N__8675\,
            I => \N__8630\
        );

    \I__2199\ : InMux
    port map (
            O => \N__8674\,
            I => \N__8625\
        );

    \I__2198\ : InMux
    port map (
            O => \N__8673\,
            I => \N__8625\
        );

    \I__2197\ : InMux
    port map (
            O => \N__8672\,
            I => \N__8622\
        );

    \I__2196\ : InMux
    port map (
            O => \N__8669\,
            I => \N__8614\
        );

    \I__2195\ : InMux
    port map (
            O => \N__8668\,
            I => \N__8614\
        );

    \I__2194\ : InMux
    port map (
            O => \N__8667\,
            I => \N__8614\
        );

    \I__2193\ : InMux
    port map (
            O => \N__8666\,
            I => \N__8609\
        );

    \I__2192\ : InMux
    port map (
            O => \N__8665\,
            I => \N__8609\
        );

    \I__2191\ : InMux
    port map (
            O => \N__8664\,
            I => \N__8604\
        );

    \I__2190\ : InMux
    port map (
            O => \N__8663\,
            I => \N__8604\
        );

    \I__2189\ : InMux
    port map (
            O => \N__8662\,
            I => \N__8601\
        );

    \I__2188\ : InMux
    port map (
            O => \N__8661\,
            I => \N__8596\
        );

    \I__2187\ : InMux
    port map (
            O => \N__8660\,
            I => \N__8596\
        );

    \I__2186\ : InMux
    port map (
            O => \N__8659\,
            I => \N__8587\
        );

    \I__2185\ : InMux
    port map (
            O => \N__8656\,
            I => \N__8587\
        );

    \I__2184\ : InMux
    port map (
            O => \N__8655\,
            I => \N__8587\
        );

    \I__2183\ : InMux
    port map (
            O => \N__8654\,
            I => \N__8587\
        );

    \I__2182\ : InMux
    port map (
            O => \N__8651\,
            I => \N__8584\
        );

    \I__2181\ : LocalMux
    port map (
            O => \N__8648\,
            I => \N__8579\
        );

    \I__2180\ : Sp12to4
    port map (
            O => \N__8645\,
            I => \N__8579\
        );

    \I__2179\ : LocalMux
    port map (
            O => \N__8642\,
            I => \N__8576\
        );

    \I__2178\ : LocalMux
    port map (
            O => \N__8639\,
            I => \N__8573\
        );

    \I__2177\ : LocalMux
    port map (
            O => \N__8636\,
            I => \N__8568\
        );

    \I__2176\ : LocalMux
    port map (
            O => \N__8633\,
            I => \N__8568\
        );

    \I__2175\ : LocalMux
    port map (
            O => \N__8630\,
            I => \N__8563\
        );

    \I__2174\ : LocalMux
    port map (
            O => \N__8625\,
            I => \N__8563\
        );

    \I__2173\ : LocalMux
    port map (
            O => \N__8622\,
            I => \N__8560\
        );

    \I__2172\ : InMux
    port map (
            O => \N__8621\,
            I => \N__8557\
        );

    \I__2171\ : LocalMux
    port map (
            O => \N__8614\,
            I => \N__8554\
        );

    \I__2170\ : LocalMux
    port map (
            O => \N__8609\,
            I => \N__8545\
        );

    \I__2169\ : LocalMux
    port map (
            O => \N__8604\,
            I => \N__8534\
        );

    \I__2168\ : LocalMux
    port map (
            O => \N__8601\,
            I => \N__8534\
        );

    \I__2167\ : LocalMux
    port map (
            O => \N__8596\,
            I => \N__8534\
        );

    \I__2166\ : LocalMux
    port map (
            O => \N__8587\,
            I => \N__8534\
        );

    \I__2165\ : LocalMux
    port map (
            O => \N__8584\,
            I => \N__8534\
        );

    \I__2164\ : Span12Mux_s3_h
    port map (
            O => \N__8579\,
            I => \N__8531\
        );

    \I__2163\ : Span4Mux_h
    port map (
            O => \N__8576\,
            I => \N__8528\
        );

    \I__2162\ : Span4Mux_h
    port map (
            O => \N__8573\,
            I => \N__8523\
        );

    \I__2161\ : Span4Mux_s3_v
    port map (
            O => \N__8568\,
            I => \N__8523\
        );

    \I__2160\ : Span4Mux_s3_v
    port map (
            O => \N__8563\,
            I => \N__8514\
        );

    \I__2159\ : Span4Mux_s3_h
    port map (
            O => \N__8560\,
            I => \N__8514\
        );

    \I__2158\ : LocalMux
    port map (
            O => \N__8557\,
            I => \N__8514\
        );

    \I__2157\ : Span4Mux_s3_h
    port map (
            O => \N__8554\,
            I => \N__8514\
        );

    \I__2156\ : InMux
    port map (
            O => \N__8553\,
            I => \N__8509\
        );

    \I__2155\ : InMux
    port map (
            O => \N__8552\,
            I => \N__8509\
        );

    \I__2154\ : InMux
    port map (
            O => \N__8551\,
            I => \N__8500\
        );

    \I__2153\ : InMux
    port map (
            O => \N__8550\,
            I => \N__8500\
        );

    \I__2152\ : InMux
    port map (
            O => \N__8549\,
            I => \N__8500\
        );

    \I__2151\ : InMux
    port map (
            O => \N__8548\,
            I => \N__8500\
        );

    \I__2150\ : Span4Mux_v
    port map (
            O => \N__8545\,
            I => \N__8495\
        );

    \I__2149\ : Span4Mux_v
    port map (
            O => \N__8534\,
            I => \N__8495\
        );

    \I__2148\ : Odrv12
    port map (
            O => \N__8531\,
            I => inc
        );

    \I__2147\ : Odrv4
    port map (
            O => \N__8528\,
            I => inc
        );

    \I__2146\ : Odrv4
    port map (
            O => \N__8523\,
            I => inc
        );

    \I__2145\ : Odrv4
    port map (
            O => \N__8514\,
            I => inc
        );

    \I__2144\ : LocalMux
    port map (
            O => \N__8509\,
            I => inc
        );

    \I__2143\ : LocalMux
    port map (
            O => \N__8500\,
            I => inc
        );

    \I__2142\ : Odrv4
    port map (
            O => \N__8495\,
            I => inc
        );

    \I__2141\ : InMux
    port map (
            O => \N__8480\,
            I => \N__8475\
        );

    \I__2140\ : InMux
    port map (
            O => \N__8479\,
            I => \N__8472\
        );

    \I__2139\ : InMux
    port map (
            O => \N__8478\,
            I => \N__8469\
        );

    \I__2138\ : LocalMux
    port map (
            O => \N__8475\,
            I => \N__8461\
        );

    \I__2137\ : LocalMux
    port map (
            O => \N__8472\,
            I => \N__8461\
        );

    \I__2136\ : LocalMux
    port map (
            O => \N__8469\,
            I => \N__8461\
        );

    \I__2135\ : InMux
    port map (
            O => \N__8468\,
            I => \N__8458\
        );

    \I__2134\ : Span4Mux_v
    port map (
            O => \N__8461\,
            I => \N__8452\
        );

    \I__2133\ : LocalMux
    port map (
            O => \N__8458\,
            I => \N__8452\
        );

    \I__2132\ : InMux
    port map (
            O => \N__8457\,
            I => \N__8449\
        );

    \I__2131\ : Span4Mux_h
    port map (
            O => \N__8452\,
            I => \N__8443\
        );

    \I__2130\ : LocalMux
    port map (
            O => \N__8449\,
            I => \N__8443\
        );

    \I__2129\ : InMux
    port map (
            O => \N__8448\,
            I => \N__8440\
        );

    \I__2128\ : Odrv4
    port map (
            O => \N__8443\,
            I => alu_out_m_0_2
        );

    \I__2127\ : LocalMux
    port map (
            O => \N__8440\,
            I => alu_out_m_0_2
        );

    \I__2126\ : InMux
    port map (
            O => \N__8435\,
            I => \N__8431\
        );

    \I__2125\ : CascadeMux
    port map (
            O => \N__8434\,
            I => \N__8428\
        );

    \I__2124\ : LocalMux
    port map (
            O => \N__8431\,
            I => \N__8422\
        );

    \I__2123\ : InMux
    port map (
            O => \N__8428\,
            I => \N__8419\
        );

    \I__2122\ : InMux
    port map (
            O => \N__8427\,
            I => \N__8416\
        );

    \I__2121\ : InMux
    port map (
            O => \N__8426\,
            I => \N__8413\
        );

    \I__2120\ : InMux
    port map (
            O => \N__8425\,
            I => \N__8408\
        );

    \I__2119\ : Span4Mux_v
    port map (
            O => \N__8422\,
            I => \N__8403\
        );

    \I__2118\ : LocalMux
    port map (
            O => \N__8419\,
            I => \N__8403\
        );

    \I__2117\ : LocalMux
    port map (
            O => \N__8416\,
            I => \N__8400\
        );

    \I__2116\ : LocalMux
    port map (
            O => \N__8413\,
            I => \N__8397\
        );

    \I__2115\ : InMux
    port map (
            O => \N__8412\,
            I => \N__8394\
        );

    \I__2114\ : InMux
    port map (
            O => \N__8411\,
            I => \N__8391\
        );

    \I__2113\ : LocalMux
    port map (
            O => \N__8408\,
            I => \N__8386\
        );

    \I__2112\ : Span4Mux_v
    port map (
            O => \N__8403\,
            I => \N__8386\
        );

    \I__2111\ : Odrv4
    port map (
            O => \N__8400\,
            I => ir_out_2
        );

    \I__2110\ : Odrv12
    port map (
            O => \N__8397\,
            I => ir_out_2
        );

    \I__2109\ : LocalMux
    port map (
            O => \N__8394\,
            I => ir_out_2
        );

    \I__2108\ : LocalMux
    port map (
            O => \N__8391\,
            I => ir_out_2
        );

    \I__2107\ : Odrv4
    port map (
            O => \N__8386\,
            I => ir_out_2
        );

    \I__2106\ : CascadeMux
    port map (
            O => \N__8375\,
            I => \N__8370\
        );

    \I__2105\ : CascadeMux
    port map (
            O => \N__8374\,
            I => \N__8365\
        );

    \I__2104\ : CascadeMux
    port map (
            O => \N__8373\,
            I => \N__8362\
        );

    \I__2103\ : InMux
    port map (
            O => \N__8370\,
            I => \N__8359\
        );

    \I__2102\ : CascadeMux
    port map (
            O => \N__8369\,
            I => \N__8356\
        );

    \I__2101\ : CascadeMux
    port map (
            O => \N__8368\,
            I => \N__8353\
        );

    \I__2100\ : InMux
    port map (
            O => \N__8365\,
            I => \N__8350\
        );

    \I__2099\ : InMux
    port map (
            O => \N__8362\,
            I => \N__8347\
        );

    \I__2098\ : LocalMux
    port map (
            O => \N__8359\,
            I => \N__8344\
        );

    \I__2097\ : InMux
    port map (
            O => \N__8356\,
            I => \N__8341\
        );

    \I__2096\ : InMux
    port map (
            O => \N__8353\,
            I => \N__8338\
        );

    \I__2095\ : LocalMux
    port map (
            O => \N__8350\,
            I => \N__8335\
        );

    \I__2094\ : LocalMux
    port map (
            O => \N__8347\,
            I => \N__8332\
        );

    \I__2093\ : Span4Mux_v
    port map (
            O => \N__8344\,
            I => \N__8325\
        );

    \I__2092\ : LocalMux
    port map (
            O => \N__8341\,
            I => \N__8325\
        );

    \I__2091\ : LocalMux
    port map (
            O => \N__8338\,
            I => \N__8325\
        );

    \I__2090\ : Span4Mux_v
    port map (
            O => \N__8335\,
            I => \N__8322\
        );

    \I__2089\ : Span4Mux_h
    port map (
            O => \N__8332\,
            I => \N__8319\
        );

    \I__2088\ : Span4Mux_h
    port map (
            O => \N__8325\,
            I => \N__8316\
        );

    \I__2087\ : Odrv4
    port map (
            O => \N__8322\,
            I => \IR_OE_2\
        );

    \I__2086\ : Odrv4
    port map (
            O => \N__8319\,
            I => \IR_OE_2\
        );

    \I__2085\ : Odrv4
    port map (
            O => \N__8316\,
            I => \IR_OE_2\
        );

    \I__2084\ : InMux
    port map (
            O => \N__8309\,
            I => \N__8303\
        );

    \I__2083\ : InMux
    port map (
            O => \N__8308\,
            I => \N__8300\
        );

    \I__2082\ : InMux
    port map (
            O => \N__8307\,
            I => \N__8297\
        );

    \I__2081\ : InMux
    port map (
            O => \N__8306\,
            I => \N__8294\
        );

    \I__2080\ : LocalMux
    port map (
            O => \N__8303\,
            I => \N__8290\
        );

    \I__2079\ : LocalMux
    port map (
            O => \N__8300\,
            I => \N__8283\
        );

    \I__2078\ : LocalMux
    port map (
            O => \N__8297\,
            I => \N__8283\
        );

    \I__2077\ : LocalMux
    port map (
            O => \N__8294\,
            I => \N__8283\
        );

    \I__2076\ : InMux
    port map (
            O => \N__8293\,
            I => \N__8280\
        );

    \I__2075\ : Span4Mux_h
    port map (
            O => \N__8290\,
            I => \N__8272\
        );

    \I__2074\ : Span4Mux_v
    port map (
            O => \N__8283\,
            I => \N__8272\
        );

    \I__2073\ : LocalMux
    port map (
            O => \N__8280\,
            I => \N__8272\
        );

    \I__2072\ : InMux
    port map (
            O => \N__8279\,
            I => \N__8269\
        );

    \I__2071\ : Span4Mux_h
    port map (
            O => \N__8272\,
            I => \N__8266\
        );

    \I__2070\ : LocalMux
    port map (
            O => \N__8269\,
            I => \N__8263\
        );

    \I__2069\ : Odrv4
    port map (
            O => \N__8266\,
            I => \pc.tbuf.g0_1_1\
        );

    \I__2068\ : Odrv4
    port map (
            O => \N__8263\,
            I => \pc.tbuf.g0_1_1\
        );

    \I__2067\ : CascadeMux
    port map (
            O => \N__8258\,
            I => \N__8254\
        );

    \I__2066\ : InMux
    port map (
            O => \N__8257\,
            I => \N__8246\
        );

    \I__2065\ : InMux
    port map (
            O => \N__8254\,
            I => \N__8246\
        );

    \I__2064\ : InMux
    port map (
            O => \N__8253\,
            I => \N__8246\
        );

    \I__2063\ : LocalMux
    port map (
            O => \N__8246\,
            I => \N__8243\
        );

    \I__2062\ : Span4Mux_h
    port map (
            O => \N__8243\,
            I => \N__8240\
        );

    \I__2061\ : Odrv4
    port map (
            O => \N__8240\,
            I => b_reg_out_2
        );

    \I__2060\ : InMux
    port map (
            O => \N__8237\,
            I => \N__8233\
        );

    \I__2059\ : InMux
    port map (
            O => \N__8236\,
            I => \N__8230\
        );

    \I__2058\ : LocalMux
    port map (
            O => \N__8233\,
            I => \N__8223\
        );

    \I__2057\ : LocalMux
    port map (
            O => \N__8230\,
            I => \N__8223\
        );

    \I__2056\ : InMux
    port map (
            O => \N__8229\,
            I => \N__8220\
        );

    \I__2055\ : InMux
    port map (
            O => \N__8228\,
            I => \N__8217\
        );

    \I__2054\ : Span4Mux_v
    port map (
            O => \N__8223\,
            I => \N__8212\
        );

    \I__2053\ : LocalMux
    port map (
            O => \N__8220\,
            I => \N__8212\
        );

    \I__2052\ : LocalMux
    port map (
            O => \N__8217\,
            I => \N__8207\
        );

    \I__2051\ : Sp12to4
    port map (
            O => \N__8212\,
            I => \N__8204\
        );

    \I__2050\ : InMux
    port map (
            O => \N__8211\,
            I => \N__8201\
        );

    \I__2049\ : InMux
    port map (
            O => \N__8210\,
            I => \N__8198\
        );

    \I__2048\ : Span12Mux_s7_v
    port map (
            O => \N__8207\,
            I => \N__8193\
        );

    \I__2047\ : Span12Mux_s8_v
    port map (
            O => \N__8204\,
            I => \N__8193\
        );

    \I__2046\ : LocalMux
    port map (
            O => \N__8201\,
            I => \N__8188\
        );

    \I__2045\ : LocalMux
    port map (
            O => \N__8198\,
            I => \N__8188\
        );

    \I__2044\ : Odrv12
    port map (
            O => \N__8193\,
            I => \IR_OE_1\
        );

    \I__2043\ : Odrv4
    port map (
            O => \N__8188\,
            I => \IR_OE_1\
        );

    \I__2042\ : InMux
    port map (
            O => \N__8183\,
            I => \N__8179\
        );

    \I__2041\ : InMux
    port map (
            O => \N__8182\,
            I => \N__8176\
        );

    \I__2040\ : LocalMux
    port map (
            O => \N__8179\,
            I => \N__8173\
        );

    \I__2039\ : LocalMux
    port map (
            O => \N__8176\,
            I => \N__8170\
        );

    \I__2038\ : Span4Mux_v
    port map (
            O => \N__8173\,
            I => \N__8161\
        );

    \I__2037\ : Span4Mux_h
    port map (
            O => \N__8170\,
            I => \N__8161\
        );

    \I__2036\ : InMux
    port map (
            O => \N__8169\,
            I => \N__8158\
        );

    \I__2035\ : InMux
    port map (
            O => \N__8168\,
            I => \N__8155\
        );

    \I__2034\ : InMux
    port map (
            O => \N__8167\,
            I => \N__8152\
        );

    \I__2033\ : InMux
    port map (
            O => \N__8166\,
            I => \N__8149\
        );

    \I__2032\ : Odrv4
    port map (
            O => \N__8161\,
            I => \pc.g0_1_0\
        );

    \I__2031\ : LocalMux
    port map (
            O => \N__8158\,
            I => \pc.g0_1_0\
        );

    \I__2030\ : LocalMux
    port map (
            O => \N__8155\,
            I => \pc.g0_1_0\
        );

    \I__2029\ : LocalMux
    port map (
            O => \N__8152\,
            I => \pc.g0_1_0\
        );

    \I__2028\ : LocalMux
    port map (
            O => \N__8149\,
            I => \pc.g0_1_0\
        );

    \I__2027\ : CascadeMux
    port map (
            O => \N__8138\,
            I => \N__8134\
        );

    \I__2026\ : CascadeMux
    port map (
            O => \N__8137\,
            I => \N__8131\
        );

    \I__2025\ : InMux
    port map (
            O => \N__8134\,
            I => \N__8126\
        );

    \I__2024\ : InMux
    port map (
            O => \N__8131\,
            I => \N__8123\
        );

    \I__2023\ : CascadeMux
    port map (
            O => \N__8130\,
            I => \N__8118\
        );

    \I__2022\ : CascadeMux
    port map (
            O => \N__8129\,
            I => \N__8115\
        );

    \I__2021\ : LocalMux
    port map (
            O => \N__8126\,
            I => \N__8109\
        );

    \I__2020\ : LocalMux
    port map (
            O => \N__8123\,
            I => \N__8109\
        );

    \I__2019\ : CascadeMux
    port map (
            O => \N__8122\,
            I => \N__8106\
        );

    \I__2018\ : CascadeMux
    port map (
            O => \N__8121\,
            I => \N__8103\
        );

    \I__2017\ : InMux
    port map (
            O => \N__8118\,
            I => \N__8100\
        );

    \I__2016\ : InMux
    port map (
            O => \N__8115\,
            I => \N__8097\
        );

    \I__2015\ : InMux
    port map (
            O => \N__8114\,
            I => \N__8094\
        );

    \I__2014\ : Span4Mux_v
    port map (
            O => \N__8109\,
            I => \N__8091\
        );

    \I__2013\ : InMux
    port map (
            O => \N__8106\,
            I => \N__8088\
        );

    \I__2012\ : InMux
    port map (
            O => \N__8103\,
            I => \N__8085\
        );

    \I__2011\ : LocalMux
    port map (
            O => \N__8100\,
            I => \N__8080\
        );

    \I__2010\ : LocalMux
    port map (
            O => \N__8097\,
            I => \N__8080\
        );

    \I__2009\ : LocalMux
    port map (
            O => \N__8094\,
            I => \N__8077\
        );

    \I__2008\ : Odrv4
    port map (
            O => \N__8091\,
            I => ir_out_1
        );

    \I__2007\ : LocalMux
    port map (
            O => \N__8088\,
            I => ir_out_1
        );

    \I__2006\ : LocalMux
    port map (
            O => \N__8085\,
            I => ir_out_1
        );

    \I__2005\ : Odrv4
    port map (
            O => \N__8080\,
            I => ir_out_1
        );

    \I__2004\ : Odrv12
    port map (
            O => \N__8077\,
            I => ir_out_1
        );

    \I__2003\ : InMux
    port map (
            O => \N__8066\,
            I => \N__8061\
        );

    \I__2002\ : InMux
    port map (
            O => \N__8065\,
            I => \N__8057\
        );

    \I__2001\ : InMux
    port map (
            O => \N__8064\,
            I => \N__8054\
        );

    \I__2000\ : LocalMux
    port map (
            O => \N__8061\,
            I => \N__8049\
        );

    \I__1999\ : InMux
    port map (
            O => \N__8060\,
            I => \N__8046\
        );

    \I__1998\ : LocalMux
    port map (
            O => \N__8057\,
            I => \N__8042\
        );

    \I__1997\ : LocalMux
    port map (
            O => \N__8054\,
            I => \N__8039\
        );

    \I__1996\ : InMux
    port map (
            O => \N__8053\,
            I => \N__8036\
        );

    \I__1995\ : InMux
    port map (
            O => \N__8052\,
            I => \N__8033\
        );

    \I__1994\ : Span4Mux_h
    port map (
            O => \N__8049\,
            I => \N__8028\
        );

    \I__1993\ : LocalMux
    port map (
            O => \N__8046\,
            I => \N__8028\
        );

    \I__1992\ : InMux
    port map (
            O => \N__8045\,
            I => \N__8025\
        );

    \I__1991\ : Odrv4
    port map (
            O => \N__8042\,
            I => alu_out_m_0_1
        );

    \I__1990\ : Odrv4
    port map (
            O => \N__8039\,
            I => alu_out_m_0_1
        );

    \I__1989\ : LocalMux
    port map (
            O => \N__8036\,
            I => alu_out_m_0_1
        );

    \I__1988\ : LocalMux
    port map (
            O => \N__8033\,
            I => alu_out_m_0_1
        );

    \I__1987\ : Odrv4
    port map (
            O => \N__8028\,
            I => alu_out_m_0_1
        );

    \I__1986\ : LocalMux
    port map (
            O => \N__8025\,
            I => alu_out_m_0_1
        );

    \I__1985\ : IoInMux
    port map (
            O => \N__8012\,
            I => \N__8009\
        );

    \I__1984\ : LocalMux
    port map (
            O => \N__8009\,
            I => \N__8006\
        );

    \I__1983\ : Odrv12
    port map (
            O => \N__8006\,
            I => out_c_1
        );

    \I__1982\ : InMux
    port map (
            O => \N__8003\,
            I => \N__7999\
        );

    \I__1981\ : InMux
    port map (
            O => \N__8002\,
            I => \N__7996\
        );

    \I__1980\ : LocalMux
    port map (
            O => \N__7999\,
            I => \N__7991\
        );

    \I__1979\ : LocalMux
    port map (
            O => \N__7996\,
            I => \N__7988\
        );

    \I__1978\ : InMux
    port map (
            O => \N__7995\,
            I => \N__7985\
        );

    \I__1977\ : InMux
    port map (
            O => \N__7994\,
            I => \N__7982\
        );

    \I__1976\ : Span4Mux_v
    port map (
            O => \N__7991\,
            I => \N__7977\
        );

    \I__1975\ : Span4Mux_h
    port map (
            O => \N__7988\,
            I => \N__7977\
        );

    \I__1974\ : LocalMux
    port map (
            O => \N__7985\,
            I => \N__7974\
        );

    \I__1973\ : LocalMux
    port map (
            O => \N__7982\,
            I => \N__7971\
        );

    \I__1972\ : Odrv4
    port map (
            O => \N__7977\,
            I => alu_out_m_4
        );

    \I__1971\ : Odrv12
    port map (
            O => \N__7974\,
            I => alu_out_m_4
        );

    \I__1970\ : Odrv4
    port map (
            O => \N__7971\,
            I => alu_out_m_4
        );

    \I__1969\ : InMux
    port map (
            O => \N__7964\,
            I => \N__7961\
        );

    \I__1968\ : LocalMux
    port map (
            O => \N__7961\,
            I => \N__7956\
        );

    \I__1967\ : InMux
    port map (
            O => \N__7960\,
            I => \N__7953\
        );

    \I__1966\ : InMux
    port map (
            O => \N__7959\,
            I => \N__7948\
        );

    \I__1965\ : Span12Mux_s3_v
    port map (
            O => \N__7956\,
            I => \N__7945\
        );

    \I__1964\ : LocalMux
    port map (
            O => \N__7953\,
            I => \N__7942\
        );

    \I__1963\ : InMux
    port map (
            O => \N__7952\,
            I => \N__7939\
        );

    \I__1962\ : InMux
    port map (
            O => \N__7951\,
            I => \N__7936\
        );

    \I__1961\ : LocalMux
    port map (
            O => \N__7948\,
            I => \N__7933\
        );

    \I__1960\ : Odrv12
    port map (
            O => \N__7945\,
            I => \mem_data_2_7_0__i2_mux_i_m\
        );

    \I__1959\ : Odrv4
    port map (
            O => \N__7942\,
            I => \mem_data_2_7_0__i2_mux_i_m\
        );

    \I__1958\ : LocalMux
    port map (
            O => \N__7939\,
            I => \mem_data_2_7_0__i2_mux_i_m\
        );

    \I__1957\ : LocalMux
    port map (
            O => \N__7936\,
            I => \mem_data_2_7_0__i2_mux_i_m\
        );

    \I__1956\ : Odrv4
    port map (
            O => \N__7933\,
            I => \mem_data_2_7_0__i2_mux_i_m\
        );

    \I__1955\ : CascadeMux
    port map (
            O => \N__7922\,
            I => \N__7919\
        );

    \I__1954\ : InMux
    port map (
            O => \N__7919\,
            I => \N__7916\
        );

    \I__1953\ : LocalMux
    port map (
            O => \N__7916\,
            I => \N__7911\
        );

    \I__1952\ : CascadeMux
    port map (
            O => \N__7915\,
            I => \N__7905\
        );

    \I__1951\ : CascadeMux
    port map (
            O => \N__7914\,
            I => \N__7900\
        );

    \I__1950\ : Span4Mux_s2_v
    port map (
            O => \N__7911\,
            I => \N__7897\
        );

    \I__1949\ : InMux
    port map (
            O => \N__7910\,
            I => \N__7892\
        );

    \I__1948\ : InMux
    port map (
            O => \N__7909\,
            I => \N__7892\
        );

    \I__1947\ : CascadeMux
    port map (
            O => \N__7908\,
            I => \N__7889\
        );

    \I__1946\ : InMux
    port map (
            O => \N__7905\,
            I => \N__7886\
        );

    \I__1945\ : CascadeMux
    port map (
            O => \N__7904\,
            I => \N__7883\
        );

    \I__1944\ : InMux
    port map (
            O => \N__7903\,
            I => \N__7878\
        );

    \I__1943\ : InMux
    port map (
            O => \N__7900\,
            I => \N__7878\
        );

    \I__1942\ : Span4Mux_h
    port map (
            O => \N__7897\,
            I => \N__7873\
        );

    \I__1941\ : LocalMux
    port map (
            O => \N__7892\,
            I => \N__7873\
        );

    \I__1940\ : InMux
    port map (
            O => \N__7889\,
            I => \N__7870\
        );

    \I__1939\ : LocalMux
    port map (
            O => \N__7886\,
            I => \N__7867\
        );

    \I__1938\ : InMux
    port map (
            O => \N__7883\,
            I => \N__7864\
        );

    \I__1937\ : LocalMux
    port map (
            O => \N__7878\,
            I => \N__7857\
        );

    \I__1936\ : Span4Mux_s2_v
    port map (
            O => \N__7873\,
            I => \N__7857\
        );

    \I__1935\ : LocalMux
    port map (
            O => \N__7870\,
            I => \N__7857\
        );

    \I__1934\ : Span4Mux_v
    port map (
            O => \N__7867\,
            I => \N__7854\
        );

    \I__1933\ : LocalMux
    port map (
            O => \N__7864\,
            I => \N__7849\
        );

    \I__1932\ : Span4Mux_v
    port map (
            O => \N__7857\,
            I => \N__7849\
        );

    \I__1931\ : Odrv4
    port map (
            O => \N__7854\,
            I => acc_out_4
        );

    \I__1930\ : Odrv4
    port map (
            O => \N__7849\,
            I => acc_out_4
        );

    \I__1929\ : IoInMux
    port map (
            O => \N__7844\,
            I => \N__7841\
        );

    \I__1928\ : LocalMux
    port map (
            O => \N__7841\,
            I => \N__7838\
        );

    \I__1927\ : Odrv12
    port map (
            O => \N__7838\,
            I => out_c_4
        );

    \I__1926\ : InMux
    port map (
            O => \N__7835\,
            I => \N__7830\
        );

    \I__1925\ : InMux
    port map (
            O => \N__7834\,
            I => \N__7825\
        );

    \I__1924\ : InMux
    port map (
            O => \N__7833\,
            I => \N__7825\
        );

    \I__1923\ : LocalMux
    port map (
            O => \N__7830\,
            I => \N__7822\
        );

    \I__1922\ : LocalMux
    port map (
            O => \N__7825\,
            I => \N__7819\
        );

    \I__1921\ : Span4Mux_h
    port map (
            O => \N__7822\,
            I => \N__7816\
        );

    \I__1920\ : Odrv4
    port map (
            O => \N__7819\,
            I => b_reg_out_3
        );

    \I__1919\ : Odrv4
    port map (
            O => \N__7816\,
            I => b_reg_out_3
        );

    \I__1918\ : CEMux
    port map (
            O => \N__7811\,
            I => \N__7808\
        );

    \I__1917\ : LocalMux
    port map (
            O => \N__7808\,
            I => \N__7805\
        );

    \I__1916\ : Span4Mux_h
    port map (
            O => \N__7805\,
            I => \N__7800\
        );

    \I__1915\ : CEMux
    port map (
            O => \N__7804\,
            I => \N__7797\
        );

    \I__1914\ : CEMux
    port map (
            O => \N__7803\,
            I => \N__7794\
        );

    \I__1913\ : Span4Mux_s2_v
    port map (
            O => \N__7800\,
            I => \N__7788\
        );

    \I__1912\ : LocalMux
    port map (
            O => \N__7797\,
            I => \N__7788\
        );

    \I__1911\ : LocalMux
    port map (
            O => \N__7794\,
            I => \N__7785\
        );

    \I__1910\ : CEMux
    port map (
            O => \N__7793\,
            I => \N__7782\
        );

    \I__1909\ : Span4Mux_v
    port map (
            O => \N__7788\,
            I => \N__7778\
        );

    \I__1908\ : Span4Mux_v
    port map (
            O => \N__7785\,
            I => \N__7773\
        );

    \I__1907\ : LocalMux
    port map (
            O => \N__7782\,
            I => \N__7773\
        );

    \I__1906\ : CEMux
    port map (
            O => \N__7781\,
            I => \N__7770\
        );

    \I__1905\ : Span4Mux_s2_v
    port map (
            O => \N__7778\,
            I => \N__7767\
        );

    \I__1904\ : Span4Mux_h
    port map (
            O => \N__7773\,
            I => \N__7764\
        );

    \I__1903\ : LocalMux
    port map (
            O => \N__7770\,
            I => \N__7761\
        );

    \I__1902\ : Odrv4
    port map (
            O => \N__7767\,
            I => \seq_B_LD_0_i\
        );

    \I__1901\ : Odrv4
    port map (
            O => \N__7764\,
            I => \seq_B_LD_0_i\
        );

    \I__1900\ : Odrv4
    port map (
            O => \N__7761\,
            I => \seq_B_LD_0_i\
        );

    \I__1899\ : InMux
    port map (
            O => \N__7754\,
            I => \N__7751\
        );

    \I__1898\ : LocalMux
    port map (
            O => \N__7751\,
            I => \N__7745\
        );

    \I__1897\ : InMux
    port map (
            O => \N__7750\,
            I => \N__7742\
        );

    \I__1896\ : InMux
    port map (
            O => \N__7749\,
            I => \N__7737\
        );

    \I__1895\ : InMux
    port map (
            O => \N__7748\,
            I => \N__7734\
        );

    \I__1894\ : Span4Mux_v
    port map (
            O => \N__7745\,
            I => \N__7729\
        );

    \I__1893\ : LocalMux
    port map (
            O => \N__7742\,
            I => \N__7729\
        );

    \I__1892\ : InMux
    port map (
            O => \N__7741\,
            I => \N__7726\
        );

    \I__1891\ : InMux
    port map (
            O => \N__7740\,
            I => \N__7723\
        );

    \I__1890\ : LocalMux
    port map (
            O => \N__7737\,
            I => \N__7720\
        );

    \I__1889\ : LocalMux
    port map (
            O => \N__7734\,
            I => \N__7717\
        );

    \I__1888\ : Span4Mux_v
    port map (
            O => \N__7729\,
            I => \N__7714\
        );

    \I__1887\ : LocalMux
    port map (
            O => \N__7726\,
            I => \N__7711\
        );

    \I__1886\ : LocalMux
    port map (
            O => \N__7723\,
            I => \N__7706\
        );

    \I__1885\ : Span4Mux_s1_h
    port map (
            O => \N__7720\,
            I => \N__7706\
        );

    \I__1884\ : Span12Mux_v
    port map (
            O => \N__7717\,
            I => \N__7703\
        );

    \I__1883\ : Span4Mux_h
    port map (
            O => \N__7714\,
            I => \N__7700\
        );

    \I__1882\ : Span4Mux_h
    port map (
            O => \N__7711\,
            I => \N__7697\
        );

    \I__1881\ : Span4Mux_v
    port map (
            O => \N__7706\,
            I => \N__7694\
        );

    \I__1880\ : Odrv12
    port map (
            O => \N__7703\,
            I => \pc.tbuf.g0_0_0\
        );

    \I__1879\ : Odrv4
    port map (
            O => \N__7700\,
            I => \pc.tbuf.g0_0_0\
        );

    \I__1878\ : Odrv4
    port map (
            O => \N__7697\,
            I => \pc.tbuf.g0_0_0\
        );

    \I__1877\ : Odrv4
    port map (
            O => \N__7694\,
            I => \pc.tbuf.g0_0_0\
        );

    \I__1876\ : InMux
    port map (
            O => \N__7685\,
            I => \N__7682\
        );

    \I__1875\ : LocalMux
    port map (
            O => \N__7682\,
            I => \N__7675\
        );

    \I__1874\ : InMux
    port map (
            O => \N__7681\,
            I => \N__7672\
        );

    \I__1873\ : InMux
    port map (
            O => \N__7680\,
            I => \N__7669\
        );

    \I__1872\ : InMux
    port map (
            O => \N__7679\,
            I => \N__7666\
        );

    \I__1871\ : InMux
    port map (
            O => \N__7678\,
            I => \N__7663\
        );

    \I__1870\ : Span4Mux_v
    port map (
            O => \N__7675\,
            I => \N__7660\
        );

    \I__1869\ : LocalMux
    port map (
            O => \N__7672\,
            I => \N__7657\
        );

    \I__1868\ : LocalMux
    port map (
            O => \N__7669\,
            I => \N__7654\
        );

    \I__1867\ : LocalMux
    port map (
            O => \N__7666\,
            I => \N__7649\
        );

    \I__1866\ : LocalMux
    port map (
            O => \N__7663\,
            I => \N__7649\
        );

    \I__1865\ : Span4Mux_h
    port map (
            O => \N__7660\,
            I => \N__7646\
        );

    \I__1864\ : Span4Mux_v
    port map (
            O => \N__7657\,
            I => \N__7643\
        );

    \I__1863\ : Span4Mux_v
    port map (
            O => \N__7654\,
            I => \N__7638\
        );

    \I__1862\ : Span4Mux_h
    port map (
            O => \N__7649\,
            I => \N__7638\
        );

    \I__1861\ : Odrv4
    port map (
            O => \N__7646\,
            I => \pc.tbuf.g0Z0Z_3\
        );

    \I__1860\ : Odrv4
    port map (
            O => \N__7643\,
            I => \pc.tbuf.g0Z0Z_3\
        );

    \I__1859\ : Odrv4
    port map (
            O => \N__7638\,
            I => \pc.tbuf.g0Z0Z_3\
        );

    \I__1858\ : CascadeMux
    port map (
            O => \N__7631\,
            I => \N__7627\
        );

    \I__1857\ : CascadeMux
    port map (
            O => \N__7630\,
            I => \N__7624\
        );

    \I__1856\ : InMux
    port map (
            O => \N__7627\,
            I => \N__7621\
        );

    \I__1855\ : InMux
    port map (
            O => \N__7624\,
            I => \N__7615\
        );

    \I__1854\ : LocalMux
    port map (
            O => \N__7621\,
            I => \N__7612\
        );

    \I__1853\ : CascadeMux
    port map (
            O => \N__7620\,
            I => \N__7609\
        );

    \I__1852\ : CascadeMux
    port map (
            O => \N__7619\,
            I => \N__7606\
        );

    \I__1851\ : InMux
    port map (
            O => \N__7618\,
            I => \N__7603\
        );

    \I__1850\ : LocalMux
    port map (
            O => \N__7615\,
            I => \N__7600\
        );

    \I__1849\ : Span4Mux_v
    port map (
            O => \N__7612\,
            I => \N__7597\
        );

    \I__1848\ : InMux
    port map (
            O => \N__7609\,
            I => \N__7594\
        );

    \I__1847\ : InMux
    port map (
            O => \N__7606\,
            I => \N__7590\
        );

    \I__1846\ : LocalMux
    port map (
            O => \N__7603\,
            I => \N__7587\
        );

    \I__1845\ : Span4Mux_v
    port map (
            O => \N__7600\,
            I => \N__7584\
        );

    \I__1844\ : Sp12to4
    port map (
            O => \N__7597\,
            I => \N__7579\
        );

    \I__1843\ : LocalMux
    port map (
            O => \N__7594\,
            I => \N__7579\
        );

    \I__1842\ : CascadeMux
    port map (
            O => \N__7593\,
            I => \N__7576\
        );

    \I__1841\ : LocalMux
    port map (
            O => \N__7590\,
            I => \N__7573\
        );

    \I__1840\ : Span4Mux_v
    port map (
            O => \N__7587\,
            I => \N__7570\
        );

    \I__1839\ : Span4Mux_h
    port map (
            O => \N__7584\,
            I => \N__7567\
        );

    \I__1838\ : Span12Mux_s10_h
    port map (
            O => \N__7579\,
            I => \N__7564\
        );

    \I__1837\ : InMux
    port map (
            O => \N__7576\,
            I => \N__7561\
        );

    \I__1836\ : Span4Mux_v
    port map (
            O => \N__7573\,
            I => \N__7556\
        );

    \I__1835\ : Span4Mux_v
    port map (
            O => \N__7570\,
            I => \N__7556\
        );

    \I__1834\ : Odrv4
    port map (
            O => \N__7567\,
            I => \pc.tbuf.gZ0Z2\
        );

    \I__1833\ : Odrv12
    port map (
            O => \N__7564\,
            I => \pc.tbuf.gZ0Z2\
        );

    \I__1832\ : LocalMux
    port map (
            O => \N__7561\,
            I => \pc.tbuf.gZ0Z2\
        );

    \I__1831\ : Odrv4
    port map (
            O => \N__7556\,
            I => \pc.tbuf.gZ0Z2\
        );

    \I__1830\ : InMux
    port map (
            O => \N__7547\,
            I => \N__7541\
        );

    \I__1829\ : InMux
    port map (
            O => \N__7546\,
            I => \N__7537\
        );

    \I__1828\ : InMux
    port map (
            O => \N__7545\,
            I => \N__7534\
        );

    \I__1827\ : InMux
    port map (
            O => \N__7544\,
            I => \N__7531\
        );

    \I__1826\ : LocalMux
    port map (
            O => \N__7541\,
            I => \N__7528\
        );

    \I__1825\ : InMux
    port map (
            O => \N__7540\,
            I => \N__7525\
        );

    \I__1824\ : LocalMux
    port map (
            O => \N__7537\,
            I => \N__7521\
        );

    \I__1823\ : LocalMux
    port map (
            O => \N__7534\,
            I => \N__7518\
        );

    \I__1822\ : LocalMux
    port map (
            O => \N__7531\,
            I => \N__7515\
        );

    \I__1821\ : Span4Mux_v
    port map (
            O => \N__7528\,
            I => \N__7510\
        );

    \I__1820\ : LocalMux
    port map (
            O => \N__7525\,
            I => \N__7510\
        );

    \I__1819\ : InMux
    port map (
            O => \N__7524\,
            I => \N__7507\
        );

    \I__1818\ : Span4Mux_h
    port map (
            O => \N__7521\,
            I => \N__7500\
        );

    \I__1817\ : Span4Mux_s3_h
    port map (
            O => \N__7518\,
            I => \N__7500\
        );

    \I__1816\ : Span4Mux_s3_h
    port map (
            O => \N__7515\,
            I => \N__7500\
        );

    \I__1815\ : Odrv4
    port map (
            O => \N__7510\,
            I => alu_out_m_1_3
        );

    \I__1814\ : LocalMux
    port map (
            O => \N__7507\,
            I => alu_out_m_1_3
        );

    \I__1813\ : Odrv4
    port map (
            O => \N__7500\,
            I => alu_out_m_1_3
        );

    \I__1812\ : IoInMux
    port map (
            O => \N__7493\,
            I => \N__7490\
        );

    \I__1811\ : LocalMux
    port map (
            O => \N__7490\,
            I => \N__7487\
        );

    \I__1810\ : Odrv12
    port map (
            O => \N__7487\,
            I => out_c_3
        );

    \I__1809\ : CEMux
    port map (
            O => \N__7484\,
            I => \N__7481\
        );

    \I__1808\ : LocalMux
    port map (
            O => \N__7481\,
            I => \N__7470\
        );

    \I__1807\ : CEMux
    port map (
            O => \N__7480\,
            I => \N__7467\
        );

    \I__1806\ : InMux
    port map (
            O => \N__7479\,
            I => \N__7464\
        );

    \I__1805\ : CEMux
    port map (
            O => \N__7478\,
            I => \N__7461\
        );

    \I__1804\ : InMux
    port map (
            O => \N__7477\,
            I => \N__7458\
        );

    \I__1803\ : InMux
    port map (
            O => \N__7476\,
            I => \N__7451\
        );

    \I__1802\ : CEMux
    port map (
            O => \N__7475\,
            I => \N__7448\
        );

    \I__1801\ : CEMux
    port map (
            O => \N__7474\,
            I => \N__7445\
        );

    \I__1800\ : CEMux
    port map (
            O => \N__7473\,
            I => \N__7442\
        );

    \I__1799\ : Span4Mux_v
    port map (
            O => \N__7470\,
            I => \N__7438\
        );

    \I__1798\ : LocalMux
    port map (
            O => \N__7467\,
            I => \N__7435\
        );

    \I__1797\ : LocalMux
    port map (
            O => \N__7464\,
            I => \N__7432\
        );

    \I__1796\ : LocalMux
    port map (
            O => \N__7461\,
            I => \N__7427\
        );

    \I__1795\ : LocalMux
    port map (
            O => \N__7458\,
            I => \N__7427\
        );

    \I__1794\ : InMux
    port map (
            O => \N__7457\,
            I => \N__7424\
        );

    \I__1793\ : InMux
    port map (
            O => \N__7456\,
            I => \N__7419\
        );

    \I__1792\ : InMux
    port map (
            O => \N__7455\,
            I => \N__7419\
        );

    \I__1791\ : InMux
    port map (
            O => \N__7454\,
            I => \N__7416\
        );

    \I__1790\ : LocalMux
    port map (
            O => \N__7451\,
            I => \N__7413\
        );

    \I__1789\ : LocalMux
    port map (
            O => \N__7448\,
            I => \N__7409\
        );

    \I__1788\ : LocalMux
    port map (
            O => \N__7445\,
            I => \N__7404\
        );

    \I__1787\ : LocalMux
    port map (
            O => \N__7442\,
            I => \N__7404\
        );

    \I__1786\ : InMux
    port map (
            O => \N__7441\,
            I => \N__7401\
        );

    \I__1785\ : Span4Mux_h
    port map (
            O => \N__7438\,
            I => \N__7389\
        );

    \I__1784\ : Span4Mux_v
    port map (
            O => \N__7435\,
            I => \N__7389\
        );

    \I__1783\ : Span4Mux_v
    port map (
            O => \N__7432\,
            I => \N__7389\
        );

    \I__1782\ : Span4Mux_h
    port map (
            O => \N__7427\,
            I => \N__7389\
        );

    \I__1781\ : LocalMux
    port map (
            O => \N__7424\,
            I => \N__7385\
        );

    \I__1780\ : LocalMux
    port map (
            O => \N__7419\,
            I => \N__7378\
        );

    \I__1779\ : LocalMux
    port map (
            O => \N__7416\,
            I => \N__7378\
        );

    \I__1778\ : Span4Mux_v
    port map (
            O => \N__7413\,
            I => \N__7378\
        );

    \I__1777\ : InMux
    port map (
            O => \N__7412\,
            I => \N__7375\
        );

    \I__1776\ : Span4Mux_h
    port map (
            O => \N__7409\,
            I => \N__7370\
        );

    \I__1775\ : Span4Mux_v
    port map (
            O => \N__7404\,
            I => \N__7370\
        );

    \I__1774\ : LocalMux
    port map (
            O => \N__7401\,
            I => \N__7367\
        );

    \I__1773\ : InMux
    port map (
            O => \N__7400\,
            I => \N__7364\
        );

    \I__1772\ : InMux
    port map (
            O => \N__7399\,
            I => \N__7361\
        );

    \I__1771\ : InMux
    port map (
            O => \N__7398\,
            I => \N__7358\
        );

    \I__1770\ : Span4Mux_h
    port map (
            O => \N__7389\,
            I => \N__7355\
        );

    \I__1769\ : InMux
    port map (
            O => \N__7388\,
            I => \N__7352\
        );

    \I__1768\ : Span4Mux_s2_v
    port map (
            O => \N__7385\,
            I => \N__7345\
        );

    \I__1767\ : Span4Mux_v
    port map (
            O => \N__7378\,
            I => \N__7345\
        );

    \I__1766\ : LocalMux
    port map (
            O => \N__7375\,
            I => \N__7345\
        );

    \I__1765\ : Span4Mux_h
    port map (
            O => \N__7370\,
            I => \N__7340\
        );

    \I__1764\ : Span4Mux_v
    port map (
            O => \N__7367\,
            I => \N__7340\
        );

    \I__1763\ : LocalMux
    port map (
            O => \N__7364\,
            I => \N__7333\
        );

    \I__1762\ : LocalMux
    port map (
            O => \N__7361\,
            I => \N__7333\
        );

    \I__1761\ : LocalMux
    port map (
            O => \N__7358\,
            I => \N__7333\
        );

    \I__1760\ : Odrv4
    port map (
            O => \N__7355\,
            I => \OUT_LD\
        );

    \I__1759\ : LocalMux
    port map (
            O => \N__7352\,
            I => \OUT_LD\
        );

    \I__1758\ : Odrv4
    port map (
            O => \N__7345\,
            I => \OUT_LD\
        );

    \I__1757\ : Odrv4
    port map (
            O => \N__7340\,
            I => \OUT_LD\
        );

    \I__1756\ : Odrv12
    port map (
            O => \N__7333\,
            I => \OUT_LD\
        );

    \I__1755\ : SRMux
    port map (
            O => \N__7322\,
            I => \N__7214\
        );

    \I__1754\ : SRMux
    port map (
            O => \N__7321\,
            I => \N__7214\
        );

    \I__1753\ : SRMux
    port map (
            O => \N__7320\,
            I => \N__7214\
        );

    \I__1752\ : SRMux
    port map (
            O => \N__7319\,
            I => \N__7214\
        );

    \I__1751\ : SRMux
    port map (
            O => \N__7318\,
            I => \N__7214\
        );

    \I__1750\ : SRMux
    port map (
            O => \N__7317\,
            I => \N__7214\
        );

    \I__1749\ : SRMux
    port map (
            O => \N__7316\,
            I => \N__7214\
        );

    \I__1748\ : SRMux
    port map (
            O => \N__7315\,
            I => \N__7214\
        );

    \I__1747\ : SRMux
    port map (
            O => \N__7314\,
            I => \N__7214\
        );

    \I__1746\ : SRMux
    port map (
            O => \N__7313\,
            I => \N__7214\
        );

    \I__1745\ : SRMux
    port map (
            O => \N__7312\,
            I => \N__7214\
        );

    \I__1744\ : SRMux
    port map (
            O => \N__7311\,
            I => \N__7214\
        );

    \I__1743\ : SRMux
    port map (
            O => \N__7310\,
            I => \N__7214\
        );

    \I__1742\ : SRMux
    port map (
            O => \N__7309\,
            I => \N__7214\
        );

    \I__1741\ : SRMux
    port map (
            O => \N__7308\,
            I => \N__7214\
        );

    \I__1740\ : SRMux
    port map (
            O => \N__7307\,
            I => \N__7214\
        );

    \I__1739\ : SRMux
    port map (
            O => \N__7306\,
            I => \N__7214\
        );

    \I__1738\ : SRMux
    port map (
            O => \N__7305\,
            I => \N__7214\
        );

    \I__1737\ : SRMux
    port map (
            O => \N__7304\,
            I => \N__7214\
        );

    \I__1736\ : SRMux
    port map (
            O => \N__7303\,
            I => \N__7214\
        );

    \I__1735\ : SRMux
    port map (
            O => \N__7302\,
            I => \N__7214\
        );

    \I__1734\ : SRMux
    port map (
            O => \N__7301\,
            I => \N__7214\
        );

    \I__1733\ : SRMux
    port map (
            O => \N__7300\,
            I => \N__7214\
        );

    \I__1732\ : SRMux
    port map (
            O => \N__7299\,
            I => \N__7214\
        );

    \I__1731\ : SRMux
    port map (
            O => \N__7298\,
            I => \N__7214\
        );

    \I__1730\ : SRMux
    port map (
            O => \N__7297\,
            I => \N__7214\
        );

    \I__1729\ : SRMux
    port map (
            O => \N__7296\,
            I => \N__7214\
        );

    \I__1728\ : SRMux
    port map (
            O => \N__7295\,
            I => \N__7214\
        );

    \I__1727\ : SRMux
    port map (
            O => \N__7294\,
            I => \N__7214\
        );

    \I__1726\ : SRMux
    port map (
            O => \N__7293\,
            I => \N__7214\
        );

    \I__1725\ : SRMux
    port map (
            O => \N__7292\,
            I => \N__7214\
        );

    \I__1724\ : SRMux
    port map (
            O => \N__7291\,
            I => \N__7214\
        );

    \I__1723\ : SRMux
    port map (
            O => \N__7290\,
            I => \N__7214\
        );

    \I__1722\ : SRMux
    port map (
            O => \N__7289\,
            I => \N__7214\
        );

    \I__1721\ : SRMux
    port map (
            O => \N__7288\,
            I => \N__7214\
        );

    \I__1720\ : SRMux
    port map (
            O => \N__7287\,
            I => \N__7214\
        );

    \I__1719\ : GlobalMux
    port map (
            O => \N__7214\,
            I => \N__7211\
        );

    \I__1718\ : gio2CtrlBuf
    port map (
            O => \N__7211\,
            I => clr_c_g
        );

    \I__1717\ : CascadeMux
    port map (
            O => \N__7208\,
            I => \mem_data_2_7_0__N_29_mux_cascade_\
        );

    \I__1716\ : IoInMux
    port map (
            O => \N__7205\,
            I => \N__7202\
        );

    \I__1715\ : LocalMux
    port map (
            O => \N__7202\,
            I => \N__7199\
        );

    \I__1714\ : Odrv12
    port map (
            O => \N__7199\,
            I => out_c_6
        );

    \I__1713\ : CascadeMux
    port map (
            O => \N__7196\,
            I => \N__7193\
        );

    \I__1712\ : InMux
    port map (
            O => \N__7193\,
            I => \N__7187\
        );

    \I__1711\ : InMux
    port map (
            O => \N__7192\,
            I => \N__7187\
        );

    \I__1710\ : LocalMux
    port map (
            O => \N__7187\,
            I => \N__7183\
        );

    \I__1709\ : InMux
    port map (
            O => \N__7186\,
            I => \N__7180\
        );

    \I__1708\ : Span4Mux_v
    port map (
            O => \N__7183\,
            I => \N__7168\
        );

    \I__1707\ : LocalMux
    port map (
            O => \N__7180\,
            I => \N__7168\
        );

    \I__1706\ : InMux
    port map (
            O => \N__7179\,
            I => \N__7156\
        );

    \I__1705\ : InMux
    port map (
            O => \N__7178\,
            I => \N__7156\
        );

    \I__1704\ : InMux
    port map (
            O => \N__7177\,
            I => \N__7156\
        );

    \I__1703\ : InMux
    port map (
            O => \N__7176\,
            I => \N__7156\
        );

    \I__1702\ : InMux
    port map (
            O => \N__7175\,
            I => \N__7156\
        );

    \I__1701\ : InMux
    port map (
            O => \N__7174\,
            I => \N__7151\
        );

    \I__1700\ : InMux
    port map (
            O => \N__7173\,
            I => \N__7151\
        );

    \I__1699\ : Span4Mux_h
    port map (
            O => \N__7168\,
            I => \N__7148\
        );

    \I__1698\ : InMux
    port map (
            O => \N__7167\,
            I => \N__7145\
        );

    \I__1697\ : LocalMux
    port map (
            O => \N__7156\,
            I => \N__7142\
        );

    \I__1696\ : LocalMux
    port map (
            O => \N__7151\,
            I => \N__7139\
        );

    \I__1695\ : Odrv4
    port map (
            O => \N__7148\,
            I => mar_out_2
        );

    \I__1694\ : LocalMux
    port map (
            O => \N__7145\,
            I => mar_out_2
        );

    \I__1693\ : Odrv4
    port map (
            O => \N__7142\,
            I => mar_out_2
        );

    \I__1692\ : Odrv12
    port map (
            O => \N__7139\,
            I => mar_out_2
        );

    \I__1691\ : InMux
    port map (
            O => \N__7130\,
            I => \N__7122\
        );

    \I__1690\ : InMux
    port map (
            O => \N__7129\,
            I => \N__7122\
        );

    \I__1689\ : CascadeMux
    port map (
            O => \N__7128\,
            I => \N__7115\
        );

    \I__1688\ : CascadeMux
    port map (
            O => \N__7127\,
            I => \N__7110\
        );

    \I__1687\ : LocalMux
    port map (
            O => \N__7122\,
            I => \N__7105\
        );

    \I__1686\ : InMux
    port map (
            O => \N__7121\,
            I => \N__7102\
        );

    \I__1685\ : InMux
    port map (
            O => \N__7120\,
            I => \N__7099\
        );

    \I__1684\ : InMux
    port map (
            O => \N__7119\,
            I => \N__7094\
        );

    \I__1683\ : InMux
    port map (
            O => \N__7118\,
            I => \N__7094\
        );

    \I__1682\ : InMux
    port map (
            O => \N__7115\,
            I => \N__7083\
        );

    \I__1681\ : InMux
    port map (
            O => \N__7114\,
            I => \N__7083\
        );

    \I__1680\ : InMux
    port map (
            O => \N__7113\,
            I => \N__7083\
        );

    \I__1679\ : InMux
    port map (
            O => \N__7110\,
            I => \N__7083\
        );

    \I__1678\ : InMux
    port map (
            O => \N__7109\,
            I => \N__7083\
        );

    \I__1677\ : InMux
    port map (
            O => \N__7108\,
            I => \N__7080\
        );

    \I__1676\ : Span4Mux_v
    port map (
            O => \N__7105\,
            I => \N__7077\
        );

    \I__1675\ : LocalMux
    port map (
            O => \N__7102\,
            I => \N__7070\
        );

    \I__1674\ : LocalMux
    port map (
            O => \N__7099\,
            I => \N__7070\
        );

    \I__1673\ : LocalMux
    port map (
            O => \N__7094\,
            I => \N__7070\
        );

    \I__1672\ : LocalMux
    port map (
            O => \N__7083\,
            I => \N__7067\
        );

    \I__1671\ : LocalMux
    port map (
            O => \N__7080\,
            I => mar_out_1
        );

    \I__1670\ : Odrv4
    port map (
            O => \N__7077\,
            I => mar_out_1
        );

    \I__1669\ : Odrv12
    port map (
            O => \N__7070\,
            I => mar_out_1
        );

    \I__1668\ : Odrv4
    port map (
            O => \N__7067\,
            I => mar_out_1
        );

    \I__1667\ : CascadeMux
    port map (
            O => \N__7058\,
            I => \N__7054\
        );

    \I__1666\ : InMux
    port map (
            O => \N__7057\,
            I => \N__7048\
        );

    \I__1665\ : InMux
    port map (
            O => \N__7054\,
            I => \N__7048\
        );

    \I__1664\ : CascadeMux
    port map (
            O => \N__7053\,
            I => \N__7039\
        );

    \I__1663\ : LocalMux
    port map (
            O => \N__7048\,
            I => \N__7036\
        );

    \I__1662\ : CascadeMux
    port map (
            O => \N__7047\,
            I => \N__7033\
        );

    \I__1661\ : CascadeMux
    port map (
            O => \N__7046\,
            I => \N__7030\
        );

    \I__1660\ : CascadeMux
    port map (
            O => \N__7045\,
            I => \N__7025\
        );

    \I__1659\ : InMux
    port map (
            O => \N__7044\,
            I => \N__7022\
        );

    \I__1658\ : CascadeMux
    port map (
            O => \N__7043\,
            I => \N__7019\
        );

    \I__1657\ : CascadeMux
    port map (
            O => \N__7042\,
            I => \N__7015\
        );

    \I__1656\ : InMux
    port map (
            O => \N__7039\,
            I => \N__7012\
        );

    \I__1655\ : Span4Mux_h
    port map (
            O => \N__7036\,
            I => \N__7009\
        );

    \I__1654\ : InMux
    port map (
            O => \N__7033\,
            I => \N__6998\
        );

    \I__1653\ : InMux
    port map (
            O => \N__7030\,
            I => \N__6998\
        );

    \I__1652\ : InMux
    port map (
            O => \N__7029\,
            I => \N__6998\
        );

    \I__1651\ : InMux
    port map (
            O => \N__7028\,
            I => \N__6998\
        );

    \I__1650\ : InMux
    port map (
            O => \N__7025\,
            I => \N__6998\
        );

    \I__1649\ : LocalMux
    port map (
            O => \N__7022\,
            I => \N__6995\
        );

    \I__1648\ : InMux
    port map (
            O => \N__7019\,
            I => \N__6988\
        );

    \I__1647\ : InMux
    port map (
            O => \N__7018\,
            I => \N__6988\
        );

    \I__1646\ : InMux
    port map (
            O => \N__7015\,
            I => \N__6988\
        );

    \I__1645\ : LocalMux
    port map (
            O => \N__7012\,
            I => \N__6985\
        );

    \I__1644\ : Span4Mux_h
    port map (
            O => \N__7009\,
            I => \N__6980\
        );

    \I__1643\ : LocalMux
    port map (
            O => \N__6998\,
            I => \N__6980\
        );

    \I__1642\ : Span12Mux_s10_v
    port map (
            O => \N__6995\,
            I => \N__6975\
        );

    \I__1641\ : LocalMux
    port map (
            O => \N__6988\,
            I => \N__6975\
        );

    \I__1640\ : Odrv4
    port map (
            O => \N__6985\,
            I => mar_out_3
        );

    \I__1639\ : Odrv4
    port map (
            O => \N__6980\,
            I => mar_out_3
        );

    \I__1638\ : Odrv12
    port map (
            O => \N__6975\,
            I => mar_out_3
        );

    \I__1637\ : InMux
    port map (
            O => \N__6968\,
            I => \N__6957\
        );

    \I__1636\ : InMux
    port map (
            O => \N__6967\,
            I => \N__6952\
        );

    \I__1635\ : InMux
    port map (
            O => \N__6966\,
            I => \N__6952\
        );

    \I__1634\ : InMux
    port map (
            O => \N__6965\,
            I => \N__6949\
        );

    \I__1633\ : InMux
    port map (
            O => \N__6964\,
            I => \N__6938\
        );

    \I__1632\ : InMux
    port map (
            O => \N__6963\,
            I => \N__6938\
        );

    \I__1631\ : InMux
    port map (
            O => \N__6962\,
            I => \N__6938\
        );

    \I__1630\ : InMux
    port map (
            O => \N__6961\,
            I => \N__6938\
        );

    \I__1629\ : InMux
    port map (
            O => \N__6960\,
            I => \N__6938\
        );

    \I__1628\ : LocalMux
    port map (
            O => \N__6957\,
            I => \N__6935\
        );

    \I__1627\ : LocalMux
    port map (
            O => \N__6952\,
            I => \N__6927\
        );

    \I__1626\ : LocalMux
    port map (
            O => \N__6949\,
            I => \N__6927\
        );

    \I__1625\ : LocalMux
    port map (
            O => \N__6938\,
            I => \N__6924\
        );

    \I__1624\ : Span4Mux_v
    port map (
            O => \N__6935\,
            I => \N__6921\
        );

    \I__1623\ : InMux
    port map (
            O => \N__6934\,
            I => \N__6914\
        );

    \I__1622\ : InMux
    port map (
            O => \N__6933\,
            I => \N__6914\
        );

    \I__1621\ : InMux
    port map (
            O => \N__6932\,
            I => \N__6914\
        );

    \I__1620\ : Span4Mux_v
    port map (
            O => \N__6927\,
            I => \N__6909\
        );

    \I__1619\ : Span4Mux_h
    port map (
            O => \N__6924\,
            I => \N__6909\
        );

    \I__1618\ : Odrv4
    port map (
            O => \N__6921\,
            I => mar_out_0
        );

    \I__1617\ : LocalMux
    port map (
            O => \N__6914\,
            I => mar_out_0
        );

    \I__1616\ : Odrv4
    port map (
            O => \N__6909\,
            I => mar_out_0
        );

    \I__1615\ : InMux
    port map (
            O => \N__6902\,
            I => \N__6895\
        );

    \I__1614\ : InMux
    port map (
            O => \N__6901\,
            I => \N__6895\
        );

    \I__1613\ : InMux
    port map (
            O => \N__6900\,
            I => \N__6892\
        );

    \I__1612\ : LocalMux
    port map (
            O => \N__6895\,
            I => \N__6887\
        );

    \I__1611\ : LocalMux
    port map (
            O => \N__6892\,
            I => \N__6884\
        );

    \I__1610\ : CascadeMux
    port map (
            O => \N__6891\,
            I => \N__6881\
        );

    \I__1609\ : CascadeMux
    port map (
            O => \N__6890\,
            I => \N__6878\
        );

    \I__1608\ : Span4Mux_s2_h
    port map (
            O => \N__6887\,
            I => \N__6875\
        );

    \I__1607\ : Span4Mux_h
    port map (
            O => \N__6884\,
            I => \N__6872\
        );

    \I__1606\ : InMux
    port map (
            O => \N__6881\,
            I => \N__6869\
        );

    \I__1605\ : InMux
    port map (
            O => \N__6878\,
            I => \N__6866\
        );

    \I__1604\ : Span4Mux_h
    port map (
            O => \N__6875\,
            I => \N__6863\
        );

    \I__1603\ : Odrv4
    port map (
            O => \N__6872\,
            I => \mem_data_2_7_0__i2_mux_0\
        );

    \I__1602\ : LocalMux
    port map (
            O => \N__6869\,
            I => \mem_data_2_7_0__i2_mux_0\
        );

    \I__1601\ : LocalMux
    port map (
            O => \N__6866\,
            I => \mem_data_2_7_0__i2_mux_0\
        );

    \I__1600\ : Odrv4
    port map (
            O => \N__6863\,
            I => \mem_data_2_7_0__i2_mux_0\
        );

    \I__1599\ : InMux
    port map (
            O => \N__6854\,
            I => \N__6851\
        );

    \I__1598\ : LocalMux
    port map (
            O => \N__6851\,
            I => \N__6848\
        );

    \I__1597\ : Span4Mux_h
    port map (
            O => \N__6848\,
            I => \N__6844\
        );

    \I__1596\ : InMux
    port map (
            O => \N__6847\,
            I => \N__6841\
        );

    \I__1595\ : Odrv4
    port map (
            O => \N__6844\,
            I => b_reg_out_1
        );

    \I__1594\ : LocalMux
    port map (
            O => \N__6841\,
            I => b_reg_out_1
        );

    \I__1593\ : CascadeMux
    port map (
            O => \N__6836\,
            I => \N__6833\
        );

    \I__1592\ : InMux
    port map (
            O => \N__6833\,
            I => \N__6830\
        );

    \I__1591\ : LocalMux
    port map (
            O => \N__6830\,
            I => \N__6826\
        );

    \I__1590\ : InMux
    port map (
            O => \N__6829\,
            I => \N__6823\
        );

    \I__1589\ : Span4Mux_s3_v
    port map (
            O => \N__6826\,
            I => \N__6817\
        );

    \I__1588\ : LocalMux
    port map (
            O => \N__6823\,
            I => \N__6814\
        );

    \I__1587\ : InMux
    port map (
            O => \N__6822\,
            I => \N__6811\
        );

    \I__1586\ : InMux
    port map (
            O => \N__6821\,
            I => \N__6808\
        );

    \I__1585\ : InMux
    port map (
            O => \N__6820\,
            I => \N__6805\
        );

    \I__1584\ : Span4Mux_s1_h
    port map (
            O => \N__6817\,
            I => \N__6800\
        );

    \I__1583\ : Span4Mux_s3_v
    port map (
            O => \N__6814\,
            I => \N__6800\
        );

    \I__1582\ : LocalMux
    port map (
            O => \N__6811\,
            I => acc_out_m_6
        );

    \I__1581\ : LocalMux
    port map (
            O => \N__6808\,
            I => acc_out_m_6
        );

    \I__1580\ : LocalMux
    port map (
            O => \N__6805\,
            I => acc_out_m_6
        );

    \I__1579\ : Odrv4
    port map (
            O => \N__6800\,
            I => acc_out_m_6
        );

    \I__1578\ : InMux
    port map (
            O => \N__6791\,
            I => \N__6786\
        );

    \I__1577\ : InMux
    port map (
            O => \N__6790\,
            I => \N__6783\
        );

    \I__1576\ : InMux
    port map (
            O => \N__6789\,
            I => \N__6779\
        );

    \I__1575\ : LocalMux
    port map (
            O => \N__6786\,
            I => \N__6775\
        );

    \I__1574\ : LocalMux
    port map (
            O => \N__6783\,
            I => \N__6772\
        );

    \I__1573\ : InMux
    port map (
            O => \N__6782\,
            I => \N__6769\
        );

    \I__1572\ : LocalMux
    port map (
            O => \N__6779\,
            I => \N__6766\
        );

    \I__1571\ : InMux
    port map (
            O => \N__6778\,
            I => \N__6763\
        );

    \I__1570\ : Span4Mux_s3_v
    port map (
            O => \N__6775\,
            I => \N__6756\
        );

    \I__1569\ : Span4Mux_s3_v
    port map (
            O => \N__6772\,
            I => \N__6756\
        );

    \I__1568\ : LocalMux
    port map (
            O => \N__6769\,
            I => \N__6756\
        );

    \I__1567\ : Span4Mux_s3_h
    port map (
            O => \N__6766\,
            I => \N__6753\
        );

    \I__1566\ : LocalMux
    port map (
            O => \N__6763\,
            I => alu_out_m_6
        );

    \I__1565\ : Odrv4
    port map (
            O => \N__6756\,
            I => alu_out_m_6
        );

    \I__1564\ : Odrv4
    port map (
            O => \N__6753\,
            I => alu_out_m_6
        );

    \I__1563\ : CascadeMux
    port map (
            O => \N__6746\,
            I => \N__6742\
        );

    \I__1562\ : InMux
    port map (
            O => \N__6745\,
            I => \N__6739\
        );

    \I__1561\ : InMux
    port map (
            O => \N__6742\,
            I => \N__6736\
        );

    \I__1560\ : LocalMux
    port map (
            O => \N__6739\,
            I => \N__6729\
        );

    \I__1559\ : LocalMux
    port map (
            O => \N__6736\,
            I => \N__6729\
        );

    \I__1558\ : CascadeMux
    port map (
            O => \N__6735\,
            I => \N__6726\
        );

    \I__1557\ : CascadeMux
    port map (
            O => \N__6734\,
            I => \N__6723\
        );

    \I__1556\ : Span4Mux_v
    port map (
            O => \N__6729\,
            I => \N__6720\
        );

    \I__1555\ : InMux
    port map (
            O => \N__6726\,
            I => \N__6717\
        );

    \I__1554\ : InMux
    port map (
            O => \N__6723\,
            I => \N__6714\
        );

    \I__1553\ : Span4Mux_h
    port map (
            O => \N__6720\,
            I => \N__6711\
        );

    \I__1552\ : LocalMux
    port map (
            O => \N__6717\,
            I => \mem_data_2_7_0__N_29_mux\
        );

    \I__1551\ : LocalMux
    port map (
            O => \N__6714\,
            I => \mem_data_2_7_0__N_29_mux\
        );

    \I__1550\ : Odrv4
    port map (
            O => \N__6711\,
            I => \mem_data_2_7_0__N_29_mux\
        );

    \I__1549\ : InMux
    port map (
            O => \N__6704\,
            I => \N__6700\
        );

    \I__1548\ : InMux
    port map (
            O => \N__6703\,
            I => \N__6697\
        );

    \I__1547\ : LocalMux
    port map (
            O => \N__6700\,
            I => b_reg_out_6
        );

    \I__1546\ : LocalMux
    port map (
            O => \N__6697\,
            I => b_reg_out_6
        );

    \I__1545\ : InMux
    port map (
            O => \N__6692\,
            I => \N__6687\
        );

    \I__1544\ : InMux
    port map (
            O => \N__6691\,
            I => \N__6684\
        );

    \I__1543\ : CascadeMux
    port map (
            O => \N__6690\,
            I => \N__6680\
        );

    \I__1542\ : LocalMux
    port map (
            O => \N__6687\,
            I => \N__6677\
        );

    \I__1541\ : LocalMux
    port map (
            O => \N__6684\,
            I => \N__6674\
        );

    \I__1540\ : InMux
    port map (
            O => \N__6683\,
            I => \N__6671\
        );

    \I__1539\ : InMux
    port map (
            O => \N__6680\,
            I => \N__6667\
        );

    \I__1538\ : Span4Mux_v
    port map (
            O => \N__6677\,
            I => \N__6664\
        );

    \I__1537\ : Span4Mux_s2_v
    port map (
            O => \N__6674\,
            I => \N__6661\
        );

    \I__1536\ : LocalMux
    port map (
            O => \N__6671\,
            I => \N__6658\
        );

    \I__1535\ : InMux
    port map (
            O => \N__6670\,
            I => \N__6655\
        );

    \I__1534\ : LocalMux
    port map (
            O => \N__6667\,
            I => \N__6652\
        );

    \I__1533\ : Odrv4
    port map (
            O => \N__6664\,
            I => acc_out_m_5
        );

    \I__1532\ : Odrv4
    port map (
            O => \N__6661\,
            I => acc_out_m_5
        );

    \I__1531\ : Odrv4
    port map (
            O => \N__6658\,
            I => acc_out_m_5
        );

    \I__1530\ : LocalMux
    port map (
            O => \N__6655\,
            I => acc_out_m_5
        );

    \I__1529\ : Odrv12
    port map (
            O => \N__6652\,
            I => acc_out_m_5
        );

    \I__1528\ : InMux
    port map (
            O => \N__6641\,
            I => \N__6638\
        );

    \I__1527\ : LocalMux
    port map (
            O => \N__6638\,
            I => \N__6631\
        );

    \I__1526\ : InMux
    port map (
            O => \N__6637\,
            I => \N__6628\
        );

    \I__1525\ : InMux
    port map (
            O => \N__6636\,
            I => \N__6625\
        );

    \I__1524\ : InMux
    port map (
            O => \N__6635\,
            I => \N__6622\
        );

    \I__1523\ : InMux
    port map (
            O => \N__6634\,
            I => \N__6619\
        );

    \I__1522\ : Span4Mux_h
    port map (
            O => \N__6631\,
            I => \N__6610\
        );

    \I__1521\ : LocalMux
    port map (
            O => \N__6628\,
            I => \N__6610\
        );

    \I__1520\ : LocalMux
    port map (
            O => \N__6625\,
            I => \N__6610\
        );

    \I__1519\ : LocalMux
    port map (
            O => \N__6622\,
            I => \N__6610\
        );

    \I__1518\ : LocalMux
    port map (
            O => \N__6619\,
            I => alu_out_m_5
        );

    \I__1517\ : Odrv4
    port map (
            O => \N__6610\,
            I => alu_out_m_5
        );

    \I__1516\ : CascadeMux
    port map (
            O => \N__6605\,
            I => \N__6601\
        );

    \I__1515\ : CascadeMux
    port map (
            O => \N__6604\,
            I => \N__6595\
        );

    \I__1514\ : InMux
    port map (
            O => \N__6601\,
            I => \N__6592\
        );

    \I__1513\ : InMux
    port map (
            O => \N__6600\,
            I => \N__6589\
        );

    \I__1512\ : CascadeMux
    port map (
            O => \N__6599\,
            I => \N__6586\
        );

    \I__1511\ : CascadeMux
    port map (
            O => \N__6598\,
            I => \N__6583\
        );

    \I__1510\ : InMux
    port map (
            O => \N__6595\,
            I => \N__6580\
        );

    \I__1509\ : LocalMux
    port map (
            O => \N__6592\,
            I => \N__6575\
        );

    \I__1508\ : LocalMux
    port map (
            O => \N__6589\,
            I => \N__6575\
        );

    \I__1507\ : InMux
    port map (
            O => \N__6586\,
            I => \N__6572\
        );

    \I__1506\ : InMux
    port map (
            O => \N__6583\,
            I => \N__6569\
        );

    \I__1505\ : LocalMux
    port map (
            O => \N__6580\,
            I => \N__6564\
        );

    \I__1504\ : Span4Mux_h
    port map (
            O => \N__6575\,
            I => \N__6564\
        );

    \I__1503\ : LocalMux
    port map (
            O => \N__6572\,
            I => m20
        );

    \I__1502\ : LocalMux
    port map (
            O => \N__6569\,
            I => m20
        );

    \I__1501\ : Odrv4
    port map (
            O => \N__6564\,
            I => m20
        );

    \I__1500\ : InMux
    port map (
            O => \N__6557\,
            I => \N__6548\
        );

    \I__1499\ : InMux
    port map (
            O => \N__6556\,
            I => \N__6543\
        );

    \I__1498\ : InMux
    port map (
            O => \N__6555\,
            I => \N__6543\
        );

    \I__1497\ : InMux
    port map (
            O => \N__6554\,
            I => \N__6538\
        );

    \I__1496\ : InMux
    port map (
            O => \N__6553\,
            I => \N__6538\
        );

    \I__1495\ : InMux
    port map (
            O => \N__6552\,
            I => \N__6531\
        );

    \I__1494\ : InMux
    port map (
            O => \N__6551\,
            I => \N__6528\
        );

    \I__1493\ : LocalMux
    port map (
            O => \N__6548\,
            I => \N__6514\
        );

    \I__1492\ : LocalMux
    port map (
            O => \N__6543\,
            I => \N__6514\
        );

    \I__1491\ : LocalMux
    port map (
            O => \N__6538\,
            I => \N__6514\
        );

    \I__1490\ : InMux
    port map (
            O => \N__6537\,
            I => \N__6511\
        );

    \I__1489\ : InMux
    port map (
            O => \N__6536\,
            I => \N__6504\
        );

    \I__1488\ : InMux
    port map (
            O => \N__6535\,
            I => \N__6504\
        );

    \I__1487\ : InMux
    port map (
            O => \N__6534\,
            I => \N__6504\
        );

    \I__1486\ : LocalMux
    port map (
            O => \N__6531\,
            I => \N__6499\
        );

    \I__1485\ : LocalMux
    port map (
            O => \N__6528\,
            I => \N__6499\
        );

    \I__1484\ : InMux
    port map (
            O => \N__6527\,
            I => \N__6496\
        );

    \I__1483\ : InMux
    port map (
            O => \N__6526\,
            I => \N__6489\
        );

    \I__1482\ : InMux
    port map (
            O => \N__6525\,
            I => \N__6489\
        );

    \I__1481\ : InMux
    port map (
            O => \N__6524\,
            I => \N__6489\
        );

    \I__1480\ : InMux
    port map (
            O => \N__6523\,
            I => \N__6486\
        );

    \I__1479\ : InMux
    port map (
            O => \N__6522\,
            I => \N__6483\
        );

    \I__1478\ : InMux
    port map (
            O => \N__6521\,
            I => \N__6479\
        );

    \I__1477\ : Span4Mux_v
    port map (
            O => \N__6514\,
            I => \N__6474\
        );

    \I__1476\ : LocalMux
    port map (
            O => \N__6511\,
            I => \N__6474\
        );

    \I__1475\ : LocalMux
    port map (
            O => \N__6504\,
            I => \N__6467\
        );

    \I__1474\ : Span4Mux_s2_v
    port map (
            O => \N__6499\,
            I => \N__6467\
        );

    \I__1473\ : LocalMux
    port map (
            O => \N__6496\,
            I => \N__6467\
        );

    \I__1472\ : LocalMux
    port map (
            O => \N__6489\,
            I => \N__6460\
        );

    \I__1471\ : LocalMux
    port map (
            O => \N__6486\,
            I => \N__6455\
        );

    \I__1470\ : LocalMux
    port map (
            O => \N__6483\,
            I => \N__6455\
        );

    \I__1469\ : InMux
    port map (
            O => \N__6482\,
            I => \N__6452\
        );

    \I__1468\ : LocalMux
    port map (
            O => \N__6479\,
            I => \N__6445\
        );

    \I__1467\ : Span4Mux_h
    port map (
            O => \N__6474\,
            I => \N__6445\
        );

    \I__1466\ : Span4Mux_h
    port map (
            O => \N__6467\,
            I => \N__6445\
        );

    \I__1465\ : InMux
    port map (
            O => \N__6466\,
            I => \N__6438\
        );

    \I__1464\ : InMux
    port map (
            O => \N__6465\,
            I => \N__6438\
        );

    \I__1463\ : InMux
    port map (
            O => \N__6464\,
            I => \N__6438\
        );

    \I__1462\ : InMux
    port map (
            O => \N__6463\,
            I => \N__6435\
        );

    \I__1461\ : Odrv12
    port map (
            O => \N__6460\,
            I => \ROM_OE\
        );

    \I__1460\ : Odrv4
    port map (
            O => \N__6455\,
            I => \ROM_OE\
        );

    \I__1459\ : LocalMux
    port map (
            O => \N__6452\,
            I => \ROM_OE\
        );

    \I__1458\ : Odrv4
    port map (
            O => \N__6445\,
            I => \ROM_OE\
        );

    \I__1457\ : LocalMux
    port map (
            O => \N__6438\,
            I => \ROM_OE\
        );

    \I__1456\ : LocalMux
    port map (
            O => \N__6435\,
            I => \ROM_OE\
        );

    \I__1455\ : IoInMux
    port map (
            O => \N__6422\,
            I => \N__6419\
        );

    \I__1454\ : LocalMux
    port map (
            O => \N__6419\,
            I => \N__6416\
        );

    \I__1453\ : Span4Mux_s1_v
    port map (
            O => \N__6416\,
            I => \N__6413\
        );

    \I__1452\ : Span4Mux_h
    port map (
            O => \N__6413\,
            I => \N__6410\
        );

    \I__1451\ : Odrv4
    port map (
            O => \N__6410\,
            I => out_c_5
        );

    \I__1450\ : IoInMux
    port map (
            O => \N__6407\,
            I => \N__6404\
        );

    \I__1449\ : LocalMux
    port map (
            O => \N__6404\,
            I => \N__6401\
        );

    \I__1448\ : Odrv12
    port map (
            O => \N__6401\,
            I => out_c_2
        );

    \I__1447\ : IoInMux
    port map (
            O => \N__6398\,
            I => \N__6395\
        );

    \I__1446\ : LocalMux
    port map (
            O => \N__6395\,
            I => \N__6392\
        );

    \I__1445\ : IoSpan4Mux
    port map (
            O => \N__6392\,
            I => \N__6389\
        );

    \I__1444\ : Span4Mux_s1_h
    port map (
            O => \N__6389\,
            I => \N__6386\
        );

    \I__1443\ : Odrv4
    port map (
            O => \N__6386\,
            I => out_c_0
        );

    \I__1442\ : CEMux
    port map (
            O => \N__6383\,
            I => \N__6379\
        );

    \I__1441\ : CEMux
    port map (
            O => \N__6382\,
            I => \N__6376\
        );

    \I__1440\ : LocalMux
    port map (
            O => \N__6379\,
            I => \N__6373\
        );

    \I__1439\ : LocalMux
    port map (
            O => \N__6376\,
            I => \N__6370\
        );

    \I__1438\ : Span4Mux_v
    port map (
            O => \N__6373\,
            I => \N__6365\
        );

    \I__1437\ : Span4Mux_v
    port map (
            O => \N__6370\,
            I => \N__6365\
        );

    \I__1436\ : Span4Mux_h
    port map (
            O => \N__6365\,
            I => \N__6362\
        );

    \I__1435\ : Odrv4
    port map (
            O => \N__6362\,
            I => \mar.MAR_LD_0_0\
        );

    \I__1434\ : InMux
    port map (
            O => \N__6359\,
            I => \N__6353\
        );

    \I__1433\ : InMux
    port map (
            O => \N__6358\,
            I => \N__6353\
        );

    \I__1432\ : LocalMux
    port map (
            O => \N__6353\,
            I => b_reg_out_5
        );

    \I__1431\ : InMux
    port map (
            O => \N__6350\,
            I => \N__6347\
        );

    \I__1430\ : LocalMux
    port map (
            O => \N__6347\,
            I => \N__6343\
        );

    \I__1429\ : InMux
    port map (
            O => \N__6346\,
            I => \N__6340\
        );

    \I__1428\ : Span4Mux_h
    port map (
            O => \N__6343\,
            I => \N__6335\
        );

    \I__1427\ : LocalMux
    port map (
            O => \N__6340\,
            I => \N__6335\
        );

    \I__1426\ : Span4Mux_v
    port map (
            O => \N__6335\,
            I => \N__6331\
        );

    \I__1425\ : InMux
    port map (
            O => \N__6334\,
            I => \N__6328\
        );

    \I__1424\ : Span4Mux_h
    port map (
            O => \N__6331\,
            I => \N__6324\
        );

    \I__1423\ : LocalMux
    port map (
            O => \N__6328\,
            I => \N__6321\
        );

    \I__1422\ : InMux
    port map (
            O => \N__6327\,
            I => \N__6318\
        );

    \I__1421\ : Odrv4
    port map (
            O => \N__6324\,
            I => acc_out_m_7
        );

    \I__1420\ : Odrv12
    port map (
            O => \N__6321\,
            I => acc_out_m_7
        );

    \I__1419\ : LocalMux
    port map (
            O => \N__6318\,
            I => acc_out_m_7
        );

    \I__1418\ : InMux
    port map (
            O => \N__6311\,
            I => \N__6306\
        );

    \I__1417\ : InMux
    port map (
            O => \N__6310\,
            I => \N__6303\
        );

    \I__1416\ : CascadeMux
    port map (
            O => \N__6309\,
            I => \N__6300\
        );

    \I__1415\ : LocalMux
    port map (
            O => \N__6306\,
            I => \N__6297\
        );

    \I__1414\ : LocalMux
    port map (
            O => \N__6303\,
            I => \N__6294\
        );

    \I__1413\ : InMux
    port map (
            O => \N__6300\,
            I => \N__6290\
        );

    \I__1412\ : Span4Mux_h
    port map (
            O => \N__6297\,
            I => \N__6285\
        );

    \I__1411\ : Span4Mux_v
    port map (
            O => \N__6294\,
            I => \N__6285\
        );

    \I__1410\ : InMux
    port map (
            O => \N__6293\,
            I => \N__6282\
        );

    \I__1409\ : LocalMux
    port map (
            O => \N__6290\,
            I => \N__6279\
        );

    \I__1408\ : Span4Mux_h
    port map (
            O => \N__6285\,
            I => \N__6276\
        );

    \I__1407\ : LocalMux
    port map (
            O => \N__6282\,
            I => alu_out_m_7
        );

    \I__1406\ : Odrv12
    port map (
            O => \N__6279\,
            I => alu_out_m_7
        );

    \I__1405\ : Odrv4
    port map (
            O => \N__6276\,
            I => alu_out_m_7
        );

    \I__1404\ : InMux
    port map (
            O => \N__6269\,
            I => \N__6265\
        );

    \I__1403\ : CascadeMux
    port map (
            O => \N__6268\,
            I => \N__6262\
        );

    \I__1402\ : LocalMux
    port map (
            O => \N__6265\,
            I => \N__6259\
        );

    \I__1401\ : InMux
    port map (
            O => \N__6262\,
            I => \N__6256\
        );

    \I__1400\ : Span4Mux_v
    port map (
            O => \N__6259\,
            I => \N__6251\
        );

    \I__1399\ : LocalMux
    port map (
            O => \N__6256\,
            I => \N__6251\
        );

    \I__1398\ : Span4Mux_h
    port map (
            O => \N__6251\,
            I => \N__6248\
        );

    \I__1397\ : Odrv4
    port map (
            O => \N__6248\,
            I => b_reg_out_7
        );

    \I__1396\ : InMux
    port map (
            O => \N__6245\,
            I => \N__6240\
        );

    \I__1395\ : InMux
    port map (
            O => \N__6244\,
            I => \N__6235\
        );

    \I__1394\ : InMux
    port map (
            O => \N__6243\,
            I => \N__6235\
        );

    \I__1393\ : LocalMux
    port map (
            O => \N__6240\,
            I => \N__6232\
        );

    \I__1392\ : LocalMux
    port map (
            O => \N__6235\,
            I => \N__6229\
        );

    \I__1391\ : Odrv12
    port map (
            O => \N__6232\,
            I => b_reg_out_0
        );

    \I__1390\ : Odrv4
    port map (
            O => \N__6229\,
            I => b_reg_out_0
        );

    \I__1389\ : CascadeMux
    port map (
            O => \N__6224\,
            I => \mem.i2_mux_cascade_\
        );

    \I__1388\ : InMux
    port map (
            O => \N__6221\,
            I => \N__6218\
        );

    \I__1387\ : LocalMux
    port map (
            O => \N__6218\,
            I => \N__6215\
        );

    \I__1386\ : Span4Mux_h
    port map (
            O => \N__6215\,
            I => \N__6212\
        );

    \I__1385\ : Odrv4
    port map (
            O => \N__6212\,
            I => \pc.N_7\
        );

    \I__1384\ : InMux
    port map (
            O => \N__6209\,
            I => \N__6206\
        );

    \I__1383\ : LocalMux
    port map (
            O => \N__6206\,
            I => \N__6202\
        );

    \I__1382\ : InMux
    port map (
            O => \N__6205\,
            I => \N__6199\
        );

    \I__1381\ : Odrv4
    port map (
            O => \N__6202\,
            I => b_reg_out_4
        );

    \I__1380\ : LocalMux
    port map (
            O => \N__6199\,
            I => b_reg_out_4
        );

    \I__1379\ : InMux
    port map (
            O => \N__6194\,
            I => \N__6187\
        );

    \I__1378\ : InMux
    port map (
            O => \N__6193\,
            I => \N__6183\
        );

    \I__1377\ : InMux
    port map (
            O => \N__6192\,
            I => \N__6180\
        );

    \I__1376\ : InMux
    port map (
            O => \N__6191\,
            I => \N__6175\
        );

    \I__1375\ : InMux
    port map (
            O => \N__6190\,
            I => \N__6175\
        );

    \I__1374\ : LocalMux
    port map (
            O => \N__6187\,
            I => \N__6172\
        );

    \I__1373\ : InMux
    port map (
            O => \N__6186\,
            I => \N__6169\
        );

    \I__1372\ : LocalMux
    port map (
            O => \N__6183\,
            I => \N__6153\
        );

    \I__1371\ : LocalMux
    port map (
            O => \N__6180\,
            I => \N__6148\
        );

    \I__1370\ : LocalMux
    port map (
            O => \N__6175\,
            I => \N__6148\
        );

    \I__1369\ : Span4Mux_v
    port map (
            O => \N__6172\,
            I => \N__6143\
        );

    \I__1368\ : LocalMux
    port map (
            O => \N__6169\,
            I => \N__6143\
        );

    \I__1367\ : InMux
    port map (
            O => \N__6168\,
            I => \N__6136\
        );

    \I__1366\ : InMux
    port map (
            O => \N__6167\,
            I => \N__6136\
        );

    \I__1365\ : InMux
    port map (
            O => \N__6166\,
            I => \N__6136\
        );

    \I__1364\ : InMux
    port map (
            O => \N__6165\,
            I => \N__6131\
        );

    \I__1363\ : InMux
    port map (
            O => \N__6164\,
            I => \N__6131\
        );

    \I__1362\ : InMux
    port map (
            O => \N__6163\,
            I => \N__6124\
        );

    \I__1361\ : InMux
    port map (
            O => \N__6162\,
            I => \N__6124\
        );

    \I__1360\ : InMux
    port map (
            O => \N__6161\,
            I => \N__6124\
        );

    \I__1359\ : InMux
    port map (
            O => \N__6160\,
            I => \N__6119\
        );

    \I__1358\ : InMux
    port map (
            O => \N__6159\,
            I => \N__6119\
        );

    \I__1357\ : InMux
    port map (
            O => \N__6158\,
            I => \N__6112\
        );

    \I__1356\ : InMux
    port map (
            O => \N__6157\,
            I => \N__6112\
        );

    \I__1355\ : InMux
    port map (
            O => \N__6156\,
            I => \N__6112\
        );

    \I__1354\ : Odrv12
    port map (
            O => \N__6153\,
            I => \seq_S0_0\
        );

    \I__1353\ : Odrv4
    port map (
            O => \N__6148\,
            I => \seq_S0_0\
        );

    \I__1352\ : Odrv4
    port map (
            O => \N__6143\,
            I => \seq_S0_0\
        );

    \I__1351\ : LocalMux
    port map (
            O => \N__6136\,
            I => \seq_S0_0\
        );

    \I__1350\ : LocalMux
    port map (
            O => \N__6131\,
            I => \seq_S0_0\
        );

    \I__1349\ : LocalMux
    port map (
            O => \N__6124\,
            I => \seq_S0_0\
        );

    \I__1348\ : LocalMux
    port map (
            O => \N__6119\,
            I => \seq_S0_0\
        );

    \I__1347\ : LocalMux
    port map (
            O => \N__6112\,
            I => \seq_S0_0\
        );

    \I__1346\ : CascadeMux
    port map (
            O => \N__6095\,
            I => \N__6092\
        );

    \I__1345\ : InMux
    port map (
            O => \N__6092\,
            I => \N__6089\
        );

    \I__1344\ : LocalMux
    port map (
            O => \N__6089\,
            I => \ALU_main.N_45\
        );

    \I__1343\ : InMux
    port map (
            O => \N__6086\,
            I => \N__6083\
        );

    \I__1342\ : LocalMux
    port map (
            O => \N__6083\,
            I => \N__6080\
        );

    \I__1341\ : Span4Mux_h
    port map (
            O => \N__6080\,
            I => \N__6076\
        );

    \I__1340\ : InMux
    port map (
            O => \N__6079\,
            I => \N__6073\
        );

    \I__1339\ : Odrv4
    port map (
            O => \N__6076\,
            I => bus_5
        );

    \I__1338\ : LocalMux
    port map (
            O => \N__6073\,
            I => bus_5
        );

    \I__1337\ : InMux
    port map (
            O => \N__6068\,
            I => \N__6064\
        );

    \I__1336\ : InMux
    port map (
            O => \N__6067\,
            I => \N__6061\
        );

    \I__1335\ : LocalMux
    port map (
            O => \N__6064\,
            I => \N__6055\
        );

    \I__1334\ : LocalMux
    port map (
            O => \N__6061\,
            I => \N__6055\
        );

    \I__1333\ : InMux
    port map (
            O => \N__6060\,
            I => \N__6052\
        );

    \I__1332\ : Span4Mux_v
    port map (
            O => \N__6055\,
            I => \N__6045\
        );

    \I__1331\ : LocalMux
    port map (
            O => \N__6052\,
            I => \N__6045\
        );

    \I__1330\ : InMux
    port map (
            O => \N__6051\,
            I => \N__6042\
        );

    \I__1329\ : InMux
    port map (
            O => \N__6050\,
            I => \N__6039\
        );

    \I__1328\ : Span4Mux_h
    port map (
            O => \N__6045\,
            I => \N__6036\
        );

    \I__1327\ : LocalMux
    port map (
            O => \N__6042\,
            I => acc_out_0
        );

    \I__1326\ : LocalMux
    port map (
            O => \N__6039\,
            I => acc_out_0
        );

    \I__1325\ : Odrv4
    port map (
            O => \N__6036\,
            I => acc_out_0
        );

    \I__1324\ : InMux
    port map (
            O => \N__6029\,
            I => \N__6025\
        );

    \I__1323\ : InMux
    port map (
            O => \N__6028\,
            I => \N__6021\
        );

    \I__1322\ : LocalMux
    port map (
            O => \N__6025\,
            I => \N__6018\
        );

    \I__1321\ : InMux
    port map (
            O => \N__6024\,
            I => \N__6015\
        );

    \I__1320\ : LocalMux
    port map (
            O => \N__6021\,
            I => \N__6011\
        );

    \I__1319\ : Span4Mux_v
    port map (
            O => \N__6018\,
            I => \N__6006\
        );

    \I__1318\ : LocalMux
    port map (
            O => \N__6015\,
            I => \N__6006\
        );

    \I__1317\ : InMux
    port map (
            O => \N__6014\,
            I => \N__6003\
        );

    \I__1316\ : Span4Mux_h
    port map (
            O => \N__6011\,
            I => \N__6000\
        );

    \I__1315\ : Odrv4
    port map (
            O => \N__6006\,
            I => acc_out_1
        );

    \I__1314\ : LocalMux
    port map (
            O => \N__6003\,
            I => acc_out_1
        );

    \I__1313\ : Odrv4
    port map (
            O => \N__6000\,
            I => acc_out_1
        );

    \I__1312\ : CascadeMux
    port map (
            O => \N__5993\,
            I => \N__5986\
        );

    \I__1311\ : InMux
    port map (
            O => \N__5992\,
            I => \N__5979\
        );

    \I__1310\ : InMux
    port map (
            O => \N__5991\,
            I => \N__5979\
        );

    \I__1309\ : InMux
    port map (
            O => \N__5990\,
            I => \N__5979\
        );

    \I__1308\ : InMux
    port map (
            O => \N__5989\,
            I => \N__5976\
        );

    \I__1307\ : InMux
    port map (
            O => \N__5986\,
            I => \N__5973\
        );

    \I__1306\ : LocalMux
    port map (
            O => \N__5979\,
            I => \N__5970\
        );

    \I__1305\ : LocalMux
    port map (
            O => \N__5976\,
            I => \N__5967\
        );

    \I__1304\ : LocalMux
    port map (
            O => \N__5973\,
            I => \N__5964\
        );

    \I__1303\ : Span4Mux_h
    port map (
            O => \N__5970\,
            I => \N__5961\
        );

    \I__1302\ : Span4Mux_v
    port map (
            O => \N__5967\,
            I => \N__5958\
        );

    \I__1301\ : Span4Mux_v
    port map (
            O => \N__5964\,
            I => \N__5955\
        );

    \I__1300\ : Odrv4
    port map (
            O => \N__5961\,
            I => acc_out_2
        );

    \I__1299\ : Odrv4
    port map (
            O => \N__5958\,
            I => acc_out_2
        );

    \I__1298\ : Odrv4
    port map (
            O => \N__5955\,
            I => acc_out_2
        );

    \I__1297\ : CEMux
    port map (
            O => \N__5948\,
            I => \N__5944\
        );

    \I__1296\ : CEMux
    port map (
            O => \N__5947\,
            I => \N__5941\
        );

    \I__1295\ : LocalMux
    port map (
            O => \N__5944\,
            I => \N__5938\
        );

    \I__1294\ : LocalMux
    port map (
            O => \N__5941\,
            I => \N__5935\
        );

    \I__1293\ : Span4Mux_v
    port map (
            O => \N__5938\,
            I => \N__5932\
        );

    \I__1292\ : Span4Mux_h
    port map (
            O => \N__5935\,
            I => \N__5929\
        );

    \I__1291\ : Odrv4
    port map (
            O => \N__5932\,
            I => \seq_ACC_LD_0_i\
        );

    \I__1290\ : Odrv4
    port map (
            O => \N__5929\,
            I => \seq_ACC_LD_0_i\
        );

    \I__1289\ : CascadeMux
    port map (
            O => \N__5924\,
            I => \N__5921\
        );

    \I__1288\ : InMux
    port map (
            O => \N__5921\,
            I => \N__5918\
        );

    \I__1287\ : LocalMux
    port map (
            O => \N__5918\,
            I => \N__5915\
        );

    \I__1286\ : Odrv4
    port map (
            O => \N__5915\,
            I => \ALU_main.N_47\
        );

    \I__1285\ : CascadeMux
    port map (
            O => \N__5912\,
            I => \N__5909\
        );

    \I__1284\ : InMux
    port map (
            O => \N__5909\,
            I => \N__5903\
        );

    \I__1283\ : InMux
    port map (
            O => \N__5908\,
            I => \N__5900\
        );

    \I__1282\ : InMux
    port map (
            O => \N__5907\,
            I => \N__5895\
        );

    \I__1281\ : InMux
    port map (
            O => \N__5906\,
            I => \N__5895\
        );

    \I__1280\ : LocalMux
    port map (
            O => \N__5903\,
            I => \N__5892\
        );

    \I__1279\ : LocalMux
    port map (
            O => \N__5900\,
            I => acc_out_6
        );

    \I__1278\ : LocalMux
    port map (
            O => \N__5895\,
            I => acc_out_6
        );

    \I__1277\ : Odrv4
    port map (
            O => \N__5892\,
            I => acc_out_6
        );

    \I__1276\ : InMux
    port map (
            O => \N__5885\,
            I => \N__5882\
        );

    \I__1275\ : LocalMux
    port map (
            O => \N__5882\,
            I => \N__5879\
        );

    \I__1274\ : Odrv4
    port map (
            O => \N__5879\,
            I => \ALU_main.un1_A_axb_6_l_ofxZ0\
        );

    \I__1273\ : InMux
    port map (
            O => \N__5876\,
            I => \N__5870\
        );

    \I__1272\ : InMux
    port map (
            O => \N__5875\,
            I => \N__5870\
        );

    \I__1271\ : LocalMux
    port map (
            O => \N__5870\,
            I => \N__5867\
        );

    \I__1270\ : Span4Mux_h
    port map (
            O => \N__5867\,
            I => \N__5863\
        );

    \I__1269\ : InMux
    port map (
            O => \N__5866\,
            I => \N__5860\
        );

    \I__1268\ : Odrv4
    port map (
            O => \N__5863\,
            I => acc_out_7
        );

    \I__1267\ : LocalMux
    port map (
            O => \N__5860\,
            I => acc_out_7
        );

    \I__1266\ : CascadeMux
    port map (
            O => \N__5855\,
            I => \N__5849\
        );

    \I__1265\ : InMux
    port map (
            O => \N__5854\,
            I => \N__5842\
        );

    \I__1264\ : InMux
    port map (
            O => \N__5853\,
            I => \N__5842\
        );

    \I__1263\ : InMux
    port map (
            O => \N__5852\,
            I => \N__5842\
        );

    \I__1262\ : InMux
    port map (
            O => \N__5849\,
            I => \N__5839\
        );

    \I__1261\ : LocalMux
    port map (
            O => \N__5842\,
            I => \N__5834\
        );

    \I__1260\ : LocalMux
    port map (
            O => \N__5839\,
            I => \N__5834\
        );

    \I__1259\ : Span4Mux_h
    port map (
            O => \N__5834\,
            I => \N__5831\
        );

    \I__1258\ : Odrv4
    port map (
            O => \N__5831\,
            I => acc_out_5
        );

    \I__1257\ : CascadeMux
    port map (
            O => \N__5828\,
            I => \N__5824\
        );

    \I__1256\ : InMux
    port map (
            O => \N__5827\,
            I => \N__5817\
        );

    \I__1255\ : InMux
    port map (
            O => \N__5824\,
            I => \N__5814\
        );

    \I__1254\ : InMux
    port map (
            O => \N__5823\,
            I => \N__5811\
        );

    \I__1253\ : InMux
    port map (
            O => \N__5822\,
            I => \N__5808\
        );

    \I__1252\ : InMux
    port map (
            O => \N__5821\,
            I => \N__5803\
        );

    \I__1251\ : InMux
    port map (
            O => \N__5820\,
            I => \N__5803\
        );

    \I__1250\ : LocalMux
    port map (
            O => \N__5817\,
            I => \N__5800\
        );

    \I__1249\ : LocalMux
    port map (
            O => \N__5814\,
            I => \N__5797\
        );

    \I__1248\ : LocalMux
    port map (
            O => \N__5811\,
            I => \N__5794\
        );

    \I__1247\ : LocalMux
    port map (
            O => \N__5808\,
            I => \N__5789\
        );

    \I__1246\ : LocalMux
    port map (
            O => \N__5803\,
            I => \N__5789\
        );

    \I__1245\ : Span4Mux_h
    port map (
            O => \N__5800\,
            I => \N__5784\
        );

    \I__1244\ : Span4Mux_h
    port map (
            O => \N__5797\,
            I => \N__5784\
        );

    \I__1243\ : Odrv4
    port map (
            O => \N__5794\,
            I => acc_out_3
        );

    \I__1242\ : Odrv4
    port map (
            O => \N__5789\,
            I => acc_out_3
        );

    \I__1241\ : Odrv4
    port map (
            O => \N__5784\,
            I => acc_out_3
        );

    \I__1240\ : InMux
    port map (
            O => \N__5777\,
            I => \N__5774\
        );

    \I__1239\ : LocalMux
    port map (
            O => \N__5774\,
            I => \N__5771\
        );

    \I__1238\ : Odrv4
    port map (
            O => \N__5771\,
            I => \ALU_main.un1_A_cry_3_c_RNI552PZ0Z2\
        );

    \I__1237\ : InMux
    port map (
            O => \N__5768\,
            I => \N__5764\
        );

    \I__1236\ : InMux
    port map (
            O => \N__5767\,
            I => \N__5757\
        );

    \I__1235\ : LocalMux
    port map (
            O => \N__5764\,
            I => \N__5754\
        );

    \I__1234\ : InMux
    port map (
            O => \N__5763\,
            I => \N__5749\
        );

    \I__1233\ : InMux
    port map (
            O => \N__5762\,
            I => \N__5749\
        );

    \I__1232\ : InMux
    port map (
            O => \N__5761\,
            I => \N__5743\
        );

    \I__1231\ : InMux
    port map (
            O => \N__5760\,
            I => \N__5738\
        );

    \I__1230\ : LocalMux
    port map (
            O => \N__5757\,
            I => \N__5735\
        );

    \I__1229\ : Span4Mux_v
    port map (
            O => \N__5754\,
            I => \N__5732\
        );

    \I__1228\ : LocalMux
    port map (
            O => \N__5749\,
            I => \N__5729\
        );

    \I__1227\ : InMux
    port map (
            O => \N__5748\,
            I => \N__5722\
        );

    \I__1226\ : InMux
    port map (
            O => \N__5747\,
            I => \N__5722\
        );

    \I__1225\ : InMux
    port map (
            O => \N__5746\,
            I => \N__5722\
        );

    \I__1224\ : LocalMux
    port map (
            O => \N__5743\,
            I => \N__5719\
        );

    \I__1223\ : InMux
    port map (
            O => \N__5742\,
            I => \N__5714\
        );

    \I__1222\ : InMux
    port map (
            O => \N__5741\,
            I => \N__5714\
        );

    \I__1221\ : LocalMux
    port map (
            O => \N__5738\,
            I => \N__5711\
        );

    \I__1220\ : Span4Mux_s3_v
    port map (
            O => \N__5735\,
            I => \N__5702\
        );

    \I__1219\ : Span4Mux_h
    port map (
            O => \N__5732\,
            I => \N__5702\
        );

    \I__1218\ : Span4Mux_v
    port map (
            O => \N__5729\,
            I => \N__5702\
        );

    \I__1217\ : LocalMux
    port map (
            O => \N__5722\,
            I => \N__5702\
        );

    \I__1216\ : Span4Mux_h
    port map (
            O => \N__5719\,
            I => \N__5697\
        );

    \I__1215\ : LocalMux
    port map (
            O => \N__5714\,
            I => \N__5697\
        );

    \I__1214\ : Span12Mux_s10_h
    port map (
            O => \N__5711\,
            I => \N__5694\
        );

    \I__1213\ : Span4Mux_h
    port map (
            O => \N__5702\,
            I => \N__5689\
        );

    \I__1212\ : Span4Mux_v
    port map (
            O => \N__5697\,
            I => \N__5689\
        );

    \I__1211\ : Odrv12
    port map (
            O => \N__5694\,
            I => \seq_un1_ALU_en_0\
        );

    \I__1210\ : Odrv4
    port map (
            O => \N__5689\,
            I => \seq_un1_ALU_en_0\
        );

    \I__1209\ : CascadeMux
    port map (
            O => \N__5684\,
            I => \N__5676\
        );

    \I__1208\ : InMux
    port map (
            O => \N__5683\,
            I => \N__5668\
        );

    \I__1207\ : InMux
    port map (
            O => \N__5682\,
            I => \N__5668\
        );

    \I__1206\ : InMux
    port map (
            O => \N__5681\,
            I => \N__5665\
        );

    \I__1205\ : InMux
    port map (
            O => \N__5680\,
            I => \N__5662\
        );

    \I__1204\ : InMux
    port map (
            O => \N__5679\,
            I => \N__5659\
        );

    \I__1203\ : InMux
    port map (
            O => \N__5676\,
            I => \N__5656\
        );

    \I__1202\ : InMux
    port map (
            O => \N__5675\,
            I => \N__5653\
        );

    \I__1201\ : InMux
    port map (
            O => \N__5674\,
            I => \N__5648\
        );

    \I__1200\ : InMux
    port map (
            O => \N__5673\,
            I => \N__5648\
        );

    \I__1199\ : LocalMux
    port map (
            O => \N__5668\,
            I => \N__5645\
        );

    \I__1198\ : LocalMux
    port map (
            O => \N__5665\,
            I => \N__5640\
        );

    \I__1197\ : LocalMux
    port map (
            O => \N__5662\,
            I => \N__5637\
        );

    \I__1196\ : LocalMux
    port map (
            O => \N__5659\,
            I => \N__5634\
        );

    \I__1195\ : LocalMux
    port map (
            O => \N__5656\,
            I => \N__5631\
        );

    \I__1194\ : LocalMux
    port map (
            O => \N__5653\,
            I => \N__5626\
        );

    \I__1193\ : LocalMux
    port map (
            O => \N__5648\,
            I => \N__5626\
        );

    \I__1192\ : Span4Mux_v
    port map (
            O => \N__5645\,
            I => \N__5623\
        );

    \I__1191\ : InMux
    port map (
            O => \N__5644\,
            I => \N__5618\
        );

    \I__1190\ : InMux
    port map (
            O => \N__5643\,
            I => \N__5618\
        );

    \I__1189\ : Span4Mux_v
    port map (
            O => \N__5640\,
            I => \N__5611\
        );

    \I__1188\ : Span4Mux_h
    port map (
            O => \N__5637\,
            I => \N__5611\
        );

    \I__1187\ : Span4Mux_v
    port map (
            O => \N__5634\,
            I => \N__5611\
        );

    \I__1186\ : Span4Mux_h
    port map (
            O => \N__5631\,
            I => \N__5602\
        );

    \I__1185\ : Span4Mux_h
    port map (
            O => \N__5626\,
            I => \N__5602\
        );

    \I__1184\ : Span4Mux_h
    port map (
            O => \N__5623\,
            I => \N__5602\
        );

    \I__1183\ : LocalMux
    port map (
            O => \N__5618\,
            I => \N__5602\
        );

    \I__1182\ : Odrv4
    port map (
            O => \N__5611\,
            I => \seq_S1_0\
        );

    \I__1181\ : Odrv4
    port map (
            O => \N__5602\,
            I => \seq_S1_0\
        );

    \I__1180\ : CascadeMux
    port map (
            O => \N__5597\,
            I => \alu_out_m_4_cascade_\
        );

    \I__1179\ : InMux
    port map (
            O => \N__5594\,
            I => \N__5591\
        );

    \I__1178\ : LocalMux
    port map (
            O => \N__5591\,
            I => \N__5587\
        );

    \I__1177\ : InMux
    port map (
            O => \N__5590\,
            I => \N__5584\
        );

    \I__1176\ : Span4Mux_s1_h
    port map (
            O => \N__5587\,
            I => \N__5581\
        );

    \I__1175\ : LocalMux
    port map (
            O => \N__5584\,
            I => \N__5578\
        );

    \I__1174\ : Span4Mux_h
    port map (
            O => \N__5581\,
            I => \N__5575\
        );

    \I__1173\ : Span4Mux_v
    port map (
            O => \N__5578\,
            I => \N__5572\
        );

    \I__1172\ : Odrv4
    port map (
            O => \N__5575\,
            I => bus_4
        );

    \I__1171\ : Odrv4
    port map (
            O => \N__5572\,
            I => bus_4
        );

    \I__1170\ : CascadeMux
    port map (
            O => \N__5567\,
            I => \bus_4_cascade_\
        );

    \I__1169\ : InMux
    port map (
            O => \N__5564\,
            I => \N__5558\
        );

    \I__1168\ : InMux
    port map (
            O => \N__5563\,
            I => \N__5555\
        );

    \I__1167\ : InMux
    port map (
            O => \N__5562\,
            I => \N__5550\
        );

    \I__1166\ : InMux
    port map (
            O => \N__5561\,
            I => \N__5550\
        );

    \I__1165\ : LocalMux
    port map (
            O => \N__5558\,
            I => \N__5542\
        );

    \I__1164\ : LocalMux
    port map (
            O => \N__5555\,
            I => \N__5539\
        );

    \I__1163\ : LocalMux
    port map (
            O => \N__5550\,
            I => \N__5536\
        );

    \I__1162\ : InMux
    port map (
            O => \N__5549\,
            I => \N__5531\
        );

    \I__1161\ : InMux
    port map (
            O => \N__5548\,
            I => \N__5531\
        );

    \I__1160\ : InMux
    port map (
            O => \N__5547\,
            I => \N__5526\
        );

    \I__1159\ : InMux
    port map (
            O => \N__5546\,
            I => \N__5526\
        );

    \I__1158\ : InMux
    port map (
            O => \N__5545\,
            I => \N__5523\
        );

    \I__1157\ : Odrv4
    port map (
            O => \N__5542\,
            I => ir_out_4
        );

    \I__1156\ : Odrv12
    port map (
            O => \N__5539\,
            I => ir_out_4
        );

    \I__1155\ : Odrv4
    port map (
            O => \N__5536\,
            I => ir_out_4
        );

    \I__1154\ : LocalMux
    port map (
            O => \N__5531\,
            I => ir_out_4
        );

    \I__1153\ : LocalMux
    port map (
            O => \N__5526\,
            I => ir_out_4
        );

    \I__1152\ : LocalMux
    port map (
            O => \N__5523\,
            I => ir_out_4
        );

    \I__1151\ : InMux
    port map (
            O => \N__5510\,
            I => \N__5507\
        );

    \I__1150\ : LocalMux
    port map (
            O => \N__5507\,
            I => \N_4_0\
        );

    \I__1149\ : InMux
    port map (
            O => \N__5504\,
            I => \N__5501\
        );

    \I__1148\ : LocalMux
    port map (
            O => \N__5501\,
            I => \N__5491\
        );

    \I__1147\ : InMux
    port map (
            O => \N__5500\,
            I => \N__5488\
        );

    \I__1146\ : InMux
    port map (
            O => \N__5499\,
            I => \N__5483\
        );

    \I__1145\ : InMux
    port map (
            O => \N__5498\,
            I => \N__5483\
        );

    \I__1144\ : InMux
    port map (
            O => \N__5497\,
            I => \N__5478\
        );

    \I__1143\ : InMux
    port map (
            O => \N__5496\,
            I => \N__5478\
        );

    \I__1142\ : InMux
    port map (
            O => \N__5495\,
            I => \N__5475\
        );

    \I__1141\ : InMux
    port map (
            O => \N__5494\,
            I => \N__5472\
        );

    \I__1140\ : Span4Mux_v
    port map (
            O => \N__5491\,
            I => \N__5469\
        );

    \I__1139\ : LocalMux
    port map (
            O => \N__5488\,
            I => ir_out_i_2_5
        );

    \I__1138\ : LocalMux
    port map (
            O => \N__5483\,
            I => ir_out_i_2_5
        );

    \I__1137\ : LocalMux
    port map (
            O => \N__5478\,
            I => ir_out_i_2_5
        );

    \I__1136\ : LocalMux
    port map (
            O => \N__5475\,
            I => ir_out_i_2_5
        );

    \I__1135\ : LocalMux
    port map (
            O => \N__5472\,
            I => ir_out_i_2_5
        );

    \I__1134\ : Odrv4
    port map (
            O => \N__5469\,
            I => ir_out_i_2_5
        );

    \I__1133\ : InMux
    port map (
            O => \N__5456\,
            I => \N__5452\
        );

    \I__1132\ : InMux
    port map (
            O => \N__5455\,
            I => \N__5449\
        );

    \I__1131\ : LocalMux
    port map (
            O => \N__5452\,
            I => \N__5440\
        );

    \I__1130\ : LocalMux
    port map (
            O => \N__5449\,
            I => \N__5437\
        );

    \I__1129\ : InMux
    port map (
            O => \N__5448\,
            I => \N__5430\
        );

    \I__1128\ : InMux
    port map (
            O => \N__5447\,
            I => \N__5430\
        );

    \I__1127\ : InMux
    port map (
            O => \N__5446\,
            I => \N__5430\
        );

    \I__1126\ : InMux
    port map (
            O => \N__5445\,
            I => \N__5427\
        );

    \I__1125\ : InMux
    port map (
            O => \N__5444\,
            I => \N__5422\
        );

    \I__1124\ : InMux
    port map (
            O => \N__5443\,
            I => \N__5422\
        );

    \I__1123\ : Span4Mux_h
    port map (
            O => \N__5440\,
            I => \N__5419\
        );

    \I__1122\ : Odrv12
    port map (
            O => \N__5437\,
            I => ir_out_4_rep1
        );

    \I__1121\ : LocalMux
    port map (
            O => \N__5430\,
            I => ir_out_4_rep1
        );

    \I__1120\ : LocalMux
    port map (
            O => \N__5427\,
            I => ir_out_4_rep1
        );

    \I__1119\ : LocalMux
    port map (
            O => \N__5422\,
            I => ir_out_4_rep1
        );

    \I__1118\ : Odrv4
    port map (
            O => \N__5419\,
            I => ir_out_4_rep1
        );

    \I__1117\ : InMux
    port map (
            O => \N__5408\,
            I => \N__5402\
        );

    \I__1116\ : CascadeMux
    port map (
            O => \N__5407\,
            I => \N__5399\
        );

    \I__1115\ : InMux
    port map (
            O => \N__5406\,
            I => \N__5394\
        );

    \I__1114\ : InMux
    port map (
            O => \N__5405\,
            I => \N__5391\
        );

    \I__1113\ : LocalMux
    port map (
            O => \N__5402\,
            I => \N__5388\
        );

    \I__1112\ : InMux
    port map (
            O => \N__5399\,
            I => \N__5385\
        );

    \I__1111\ : InMux
    port map (
            O => \N__5398\,
            I => \N__5380\
        );

    \I__1110\ : InMux
    port map (
            O => \N__5397\,
            I => \N__5380\
        );

    \I__1109\ : LocalMux
    port map (
            O => \N__5394\,
            I => \N__5377\
        );

    \I__1108\ : LocalMux
    port map (
            O => \N__5391\,
            I => \IR_ff7_q_0_fast\
        );

    \I__1107\ : Odrv4
    port map (
            O => \N__5388\,
            I => \IR_ff7_q_0_fast\
        );

    \I__1106\ : LocalMux
    port map (
            O => \N__5385\,
            I => \IR_ff7_q_0_fast\
        );

    \I__1105\ : LocalMux
    port map (
            O => \N__5380\,
            I => \IR_ff7_q_0_fast\
        );

    \I__1104\ : Odrv4
    port map (
            O => \N__5377\,
            I => \IR_ff7_q_0_fast\
        );

    \I__1103\ : InMux
    port map (
            O => \N__5366\,
            I => \N__5359\
        );

    \I__1102\ : InMux
    port map (
            O => \N__5365\,
            I => \N__5354\
        );

    \I__1101\ : InMux
    port map (
            O => \N__5364\,
            I => \N__5354\
        );

    \I__1100\ : InMux
    port map (
            O => \N__5363\,
            I => \N__5351\
        );

    \I__1099\ : CascadeMux
    port map (
            O => \N__5362\,
            I => \N__5347\
        );

    \I__1098\ : LocalMux
    port map (
            O => \N__5359\,
            I => \N__5342\
        );

    \I__1097\ : LocalMux
    port map (
            O => \N__5354\,
            I => \N__5342\
        );

    \I__1096\ : LocalMux
    port map (
            O => \N__5351\,
            I => \N__5339\
        );

    \I__1095\ : InMux
    port map (
            O => \N__5350\,
            I => \N__5334\
        );

    \I__1094\ : InMux
    port map (
            O => \N__5347\,
            I => \N__5334\
        );

    \I__1093\ : Span4Mux_v
    port map (
            O => \N__5342\,
            I => \N__5327\
        );

    \I__1092\ : Span4Mux_h
    port map (
            O => \N__5339\,
            I => \N__5327\
        );

    \I__1091\ : LocalMux
    port map (
            O => \N__5334\,
            I => \N__5327\
        );

    \I__1090\ : Span4Mux_h
    port map (
            O => \N__5327\,
            I => \N__5322\
        );

    \I__1089\ : InMux
    port map (
            O => \N__5326\,
            I => \N__5317\
        );

    \I__1088\ : InMux
    port map (
            O => \N__5325\,
            I => \N__5317\
        );

    \I__1087\ : Odrv4
    port map (
            O => \N__5322\,
            I => \seq.counter.TZ0Z_4\
        );

    \I__1086\ : LocalMux
    port map (
            O => \N__5317\,
            I => \seq.counter.TZ0Z_4\
        );

    \I__1085\ : InMux
    port map (
            O => \N__5312\,
            I => \N__5306\
        );

    \I__1084\ : InMux
    port map (
            O => \N__5311\,
            I => \N__5303\
        );

    \I__1083\ : InMux
    port map (
            O => \N__5310\,
            I => \N__5300\
        );

    \I__1082\ : InMux
    port map (
            O => \N__5309\,
            I => \N__5296\
        );

    \I__1081\ : LocalMux
    port map (
            O => \N__5306\,
            I => \N__5292\
        );

    \I__1080\ : LocalMux
    port map (
            O => \N__5303\,
            I => \N__5285\
        );

    \I__1079\ : LocalMux
    port map (
            O => \N__5300\,
            I => \N__5285\
        );

    \I__1078\ : CascadeMux
    port map (
            O => \N__5299\,
            I => \N__5282\
        );

    \I__1077\ : LocalMux
    port map (
            O => \N__5296\,
            I => \N__5278\
        );

    \I__1076\ : InMux
    port map (
            O => \N__5295\,
            I => \N__5275\
        );

    \I__1075\ : Span4Mux_h
    port map (
            O => \N__5292\,
            I => \N__5272\
        );

    \I__1074\ : InMux
    port map (
            O => \N__5291\,
            I => \N__5267\
        );

    \I__1073\ : InMux
    port map (
            O => \N__5290\,
            I => \N__5267\
        );

    \I__1072\ : Span4Mux_h
    port map (
            O => \N__5285\,
            I => \N__5264\
        );

    \I__1071\ : InMux
    port map (
            O => \N__5282\,
            I => \N__5259\
        );

    \I__1070\ : InMux
    port map (
            O => \N__5281\,
            I => \N__5259\
        );

    \I__1069\ : Odrv4
    port map (
            O => \N__5278\,
            I => ir_out_7
        );

    \I__1068\ : LocalMux
    port map (
            O => \N__5275\,
            I => ir_out_7
        );

    \I__1067\ : Odrv4
    port map (
            O => \N__5272\,
            I => ir_out_7
        );

    \I__1066\ : LocalMux
    port map (
            O => \N__5267\,
            I => ir_out_7
        );

    \I__1065\ : Odrv4
    port map (
            O => \N__5264\,
            I => ir_out_7
        );

    \I__1064\ : LocalMux
    port map (
            O => \N__5259\,
            I => ir_out_7
        );

    \I__1063\ : CascadeMux
    port map (
            O => \N__5246\,
            I => \seq.g0_i_a3_0Z0Z_2_cascade_\
        );

    \I__1062\ : InMux
    port map (
            O => \N__5243\,
            I => \N__5240\
        );

    \I__1061\ : LocalMux
    port map (
            O => \N__5240\,
            I => \N__5237\
        );

    \I__1060\ : Span4Mux_h
    port map (
            O => \N__5237\,
            I => \N__5234\
        );

    \I__1059\ : Odrv4
    port map (
            O => \N__5234\,
            I => \seq.g0_i_a3Z0Z_2\
        );

    \I__1058\ : CascadeMux
    port map (
            O => \N__5231\,
            I => \seq_S0_0_cascade_\
        );

    \I__1057\ : InMux
    port map (
            O => \N__5228\,
            I => \N__5225\
        );

    \I__1056\ : LocalMux
    port map (
            O => \N__5225\,
            I => \ALU_main.un1_A_axb_5_l_ofxZ0\
        );

    \I__1055\ : InMux
    port map (
            O => \N__5222\,
            I => \N__5219\
        );

    \I__1054\ : LocalMux
    port map (
            O => \N__5219\,
            I => \N__5213\
        );

    \I__1053\ : InMux
    port map (
            O => \N__5218\,
            I => \N__5210\
        );

    \I__1052\ : InMux
    port map (
            O => \N__5217\,
            I => \N__5207\
        );

    \I__1051\ : InMux
    port map (
            O => \N__5216\,
            I => \N__5204\
        );

    \I__1050\ : Span4Mux_s3_v
    port map (
            O => \N__5213\,
            I => \N__5197\
        );

    \I__1049\ : LocalMux
    port map (
            O => \N__5210\,
            I => \N__5197\
        );

    \I__1048\ : LocalMux
    port map (
            O => \N__5207\,
            I => \N__5192\
        );

    \I__1047\ : LocalMux
    port map (
            O => \N__5204\,
            I => \N__5192\
        );

    \I__1046\ : InMux
    port map (
            O => \N__5203\,
            I => \N__5189\
        );

    \I__1045\ : CascadeMux
    port map (
            O => \N__5202\,
            I => \N__5185\
        );

    \I__1044\ : Span4Mux_v
    port map (
            O => \N__5197\,
            I => \N__5182\
        );

    \I__1043\ : Span4Mux_v
    port map (
            O => \N__5192\,
            I => \N__5179\
        );

    \I__1042\ : LocalMux
    port map (
            O => \N__5189\,
            I => \N__5176\
        );

    \I__1041\ : InMux
    port map (
            O => \N__5188\,
            I => \N__5173\
        );

    \I__1040\ : InMux
    port map (
            O => \N__5185\,
            I => \N__5170\
        );

    \I__1039\ : Span4Mux_s1_h
    port map (
            O => \N__5182\,
            I => \N__5165\
        );

    \I__1038\ : Span4Mux_s1_h
    port map (
            O => \N__5179\,
            I => \N__5165\
        );

    \I__1037\ : Odrv12
    port map (
            O => \N__5176\,
            I => \seq.counter.TZ0Z_3\
        );

    \I__1036\ : LocalMux
    port map (
            O => \N__5173\,
            I => \seq.counter.TZ0Z_3\
        );

    \I__1035\ : LocalMux
    port map (
            O => \N__5170\,
            I => \seq.counter.TZ0Z_3\
        );

    \I__1034\ : Odrv4
    port map (
            O => \N__5165\,
            I => \seq.counter.TZ0Z_3\
        );

    \I__1033\ : InMux
    port map (
            O => \N__5156\,
            I => \N__5151\
        );

    \I__1032\ : InMux
    port map (
            O => \N__5155\,
            I => \N__5148\
        );

    \I__1031\ : InMux
    port map (
            O => \N__5154\,
            I => \N__5144\
        );

    \I__1030\ : LocalMux
    port map (
            O => \N__5151\,
            I => \N__5139\
        );

    \I__1029\ : LocalMux
    port map (
            O => \N__5148\,
            I => \N__5139\
        );

    \I__1028\ : CascadeMux
    port map (
            O => \N__5147\,
            I => \N__5135\
        );

    \I__1027\ : LocalMux
    port map (
            O => \N__5144\,
            I => \N__5130\
        );

    \I__1026\ : Span4Mux_h
    port map (
            O => \N__5139\,
            I => \N__5127\
        );

    \I__1025\ : InMux
    port map (
            O => \N__5138\,
            I => \N__5120\
        );

    \I__1024\ : InMux
    port map (
            O => \N__5135\,
            I => \N__5120\
        );

    \I__1023\ : InMux
    port map (
            O => \N__5134\,
            I => \N__5120\
        );

    \I__1022\ : InMux
    port map (
            O => \N__5133\,
            I => \N__5117\
        );

    \I__1021\ : Odrv12
    port map (
            O => \N__5130\,
            I => \seq.D_2\
        );

    \I__1020\ : Odrv4
    port map (
            O => \N__5127\,
            I => \seq.D_2\
        );

    \I__1019\ : LocalMux
    port map (
            O => \N__5120\,
            I => \seq.D_2\
        );

    \I__1018\ : LocalMux
    port map (
            O => \N__5117\,
            I => \seq.D_2\
        );

    \I__1017\ : CascadeMux
    port map (
            O => \N__5108\,
            I => \N__5105\
        );

    \I__1016\ : InMux
    port map (
            O => \N__5105\,
            I => \N__5102\
        );

    \I__1015\ : LocalMux
    port map (
            O => \N__5102\,
            I => \N__5099\
        );

    \I__1014\ : Odrv4
    port map (
            O => \N__5099\,
            I => \seq.B_LD_0_2_tz\
        );

    \I__1013\ : InMux
    port map (
            O => \N__5096\,
            I => \N__5093\
        );

    \I__1012\ : LocalMux
    port map (
            O => \N__5093\,
            I => \N__5089\
        );

    \I__1011\ : InMux
    port map (
            O => \N__5092\,
            I => \N__5085\
        );

    \I__1010\ : Span4Mux_v
    port map (
            O => \N__5089\,
            I => \N__5082\
        );

    \I__1009\ : InMux
    port map (
            O => \N__5088\,
            I => \N__5079\
        );

    \I__1008\ : LocalMux
    port map (
            O => \N__5085\,
            I => \N__5075\
        );

    \I__1007\ : Span4Mux_h
    port map (
            O => \N__5082\,
            I => \N__5070\
        );

    \I__1006\ : LocalMux
    port map (
            O => \N__5079\,
            I => \N__5070\
        );

    \I__1005\ : InMux
    port map (
            O => \N__5078\,
            I => \N__5067\
        );

    \I__1004\ : Odrv12
    port map (
            O => \N__5075\,
            I => \seq.D_1\
        );

    \I__1003\ : Odrv4
    port map (
            O => \N__5070\,
            I => \seq.D_1\
        );

    \I__1002\ : LocalMux
    port map (
            O => \N__5067\,
            I => \seq.D_1\
        );

    \I__1001\ : CascadeMux
    port map (
            O => \N__5060\,
            I => \N__5057\
        );

    \I__1000\ : InMux
    port map (
            O => \N__5057\,
            I => \N__5054\
        );

    \I__999\ : LocalMux
    port map (
            O => \N__5054\,
            I => \ALU_main.un1_A_axb_1_l_ofxZ0\
        );

    \I__998\ : InMux
    port map (
            O => \N__5051\,
            I => \N__5048\
        );

    \I__997\ : LocalMux
    port map (
            O => \N__5048\,
            I => \ALU_main.un1_A_axb_4_l_ofxZ0\
        );

    \I__996\ : CascadeMux
    port map (
            O => \N__5045\,
            I => \ALU_main_N_42_0_cascade_\
        );

    \I__995\ : InMux
    port map (
            O => \N__5042\,
            I => \N__5039\
        );

    \I__994\ : LocalMux
    port map (
            O => \N__5039\,
            I => \un1_A_cry_0_c_RNIPCLO2\
        );

    \I__993\ : CascadeMux
    port map (
            O => \N__5036\,
            I => \ALU_main_N_41_0_cascade_\
        );

    \I__992\ : InMux
    port map (
            O => \N__5033\,
            I => \N__5030\
        );

    \I__991\ : LocalMux
    port map (
            O => \N__5030\,
            I => \N__5026\
        );

    \I__990\ : InMux
    port map (
            O => \N__5029\,
            I => \N__5023\
        );

    \I__989\ : Span4Mux_s3_h
    port map (
            O => \N__5026\,
            I => \N__5020\
        );

    \I__988\ : LocalMux
    port map (
            O => \N__5023\,
            I => \un1_A_cry_0_s\
        );

    \I__987\ : Odrv4
    port map (
            O => \N__5020\,
            I => \un1_A_cry_0_s\
        );

    \I__986\ : InMux
    port map (
            O => \N__5015\,
            I => \N__5009\
        );

    \I__985\ : InMux
    port map (
            O => \N__5014\,
            I => \N__5009\
        );

    \I__984\ : LocalMux
    port map (
            O => \N__5009\,
            I => \N__5006\
        );

    \I__983\ : Span4Mux_h
    port map (
            O => \N__5006\,
            I => \N__4999\
        );

    \I__982\ : InMux
    port map (
            O => \N__5005\,
            I => \N__4992\
        );

    \I__981\ : InMux
    port map (
            O => \N__5004\,
            I => \N__4992\
        );

    \I__980\ : InMux
    port map (
            O => \N__5003\,
            I => \N__4992\
        );

    \I__979\ : InMux
    port map (
            O => \N__5002\,
            I => \N__4989\
        );

    \I__978\ : Odrv4
    port map (
            O => \N__4999\,
            I => \seq.D_4\
        );

    \I__977\ : LocalMux
    port map (
            O => \N__4992\,
            I => \seq.D_4\
        );

    \I__976\ : LocalMux
    port map (
            O => \N__4989\,
            I => \seq.D_4\
        );

    \I__975\ : InMux
    port map (
            O => \N__4982\,
            I => \N__4977\
        );

    \I__974\ : InMux
    port map (
            O => \N__4981\,
            I => \N__4972\
        );

    \I__973\ : InMux
    port map (
            O => \N__4980\,
            I => \N__4972\
        );

    \I__972\ : LocalMux
    port map (
            O => \N__4977\,
            I => \N__4969\
        );

    \I__971\ : LocalMux
    port map (
            O => \N__4972\,
            I => \N__4966\
        );

    \I__970\ : Span4Mux_v
    port map (
            O => \N__4969\,
            I => \N__4958\
        );

    \I__969\ : Span4Mux_v
    port map (
            O => \N__4966\,
            I => \N__4958\
        );

    \I__968\ : InMux
    port map (
            O => \N__4965\,
            I => \N__4953\
        );

    \I__967\ : InMux
    port map (
            O => \N__4964\,
            I => \N__4953\
        );

    \I__966\ : InMux
    port map (
            O => \N__4963\,
            I => \N__4950\
        );

    \I__965\ : Odrv4
    port map (
            O => \N__4958\,
            I => \seq.DZ0Z_0\
        );

    \I__964\ : LocalMux
    port map (
            O => \N__4953\,
            I => \seq.DZ0Z_0\
        );

    \I__963\ : LocalMux
    port map (
            O => \N__4950\,
            I => \seq.DZ0Z_0\
        );

    \I__962\ : CascadeMux
    port map (
            O => \N__4943\,
            I => \N__4940\
        );

    \I__961\ : InMux
    port map (
            O => \N__4940\,
            I => \N__4937\
        );

    \I__960\ : LocalMux
    port map (
            O => \N__4937\,
            I => \N__4934\
        );

    \I__959\ : Span4Mux_h
    port map (
            O => \N__4934\,
            I => \N__4931\
        );

    \I__958\ : Odrv4
    port map (
            O => \N__4931\,
            I => \seq.g2Z0Z_1\
        );

    \I__957\ : CascadeMux
    port map (
            O => \N__4928\,
            I => \N__4925\
        );

    \I__956\ : InMux
    port map (
            O => \N__4925\,
            I => \N__4922\
        );

    \I__955\ : LocalMux
    port map (
            O => \N__4922\,
            I => \ALU_main.un1_A_axb_0_l_ofxZ0\
        );

    \I__954\ : InMux
    port map (
            O => \N__4919\,
            I => \N__4916\
        );

    \I__953\ : LocalMux
    port map (
            O => \N__4916\,
            I => \ALU_main.un1_A_axb_3_l_ofxZ0\
        );

    \I__952\ : InMux
    port map (
            O => \N__4913\,
            I => \N__4910\
        );

    \I__951\ : LocalMux
    port map (
            O => \N__4910\,
            I => \ALU_main.un1_A_cry_4_c_RNI9D6PZ0Z2\
        );

    \I__950\ : CascadeMux
    port map (
            O => \N__4907\,
            I => \ALU_main.N_46_cascade_\
        );

    \I__949\ : InMux
    port map (
            O => \N__4904\,
            I => \N__4901\
        );

    \I__948\ : LocalMux
    port map (
            O => \N__4901\,
            I => \N__4898\
        );

    \I__947\ : Span4Mux_v
    port map (
            O => \N__4898\,
            I => \N__4894\
        );

    \I__946\ : InMux
    port map (
            O => \N__4897\,
            I => \N__4891\
        );

    \I__945\ : Span4Mux_h
    port map (
            O => \N__4894\,
            I => \N__4884\
        );

    \I__944\ : LocalMux
    port map (
            O => \N__4891\,
            I => \N__4884\
        );

    \I__943\ : InMux
    port map (
            O => \N__4890\,
            I => \N__4879\
        );

    \I__942\ : InMux
    port map (
            O => \N__4889\,
            I => \N__4879\
        );

    \I__941\ : Odrv4
    port map (
            O => \N__4884\,
            I => \seq.D_3\
        );

    \I__940\ : LocalMux
    port map (
            O => \N__4879\,
            I => \seq.D_3\
        );

    \I__939\ : CascadeMux
    port map (
            O => \N__4874\,
            I => \seq.counter.ACC_LD_0_0_cascade_\
        );

    \I__938\ : InMux
    port map (
            O => \N__4871\,
            I => \N__4868\
        );

    \I__937\ : LocalMux
    port map (
            O => \N__4868\,
            I => \N__4865\
        );

    \I__936\ : Odrv12
    port map (
            O => \N__4865\,
            I => \pc.program_counter_m_0_1\
        );

    \I__935\ : InMux
    port map (
            O => \N__4862\,
            I => \N__4859\
        );

    \I__934\ : LocalMux
    port map (
            O => \N__4859\,
            I => \pc.tbuf.out_1_1_ivZ0Z_0\
        );

    \I__933\ : CascadeMux
    port map (
            O => \N__4856\,
            I => \mem_data_2_7_0__N_11_0_cascade_\
        );

    \I__932\ : InMux
    port map (
            O => \N__4853\,
            I => \N__4850\
        );

    \I__931\ : LocalMux
    port map (
            O => \N__4850\,
            I => \pc.program_counter_4_rn_2_1\
        );

    \I__930\ : InMux
    port map (
            O => \N__4847\,
            I => \N__4844\
        );

    \I__929\ : LocalMux
    port map (
            O => \N__4844\,
            I => \pc.program_counter_4_sn_1\
        );

    \I__928\ : CascadeMux
    port map (
            O => \N__4841\,
            I => \pc.g0_1_0_cascade_\
        );

    \I__927\ : CascadeMux
    port map (
            O => \N__4838\,
            I => \N__4834\
        );

    \I__926\ : InMux
    port map (
            O => \N__4837\,
            I => \N__4829\
        );

    \I__925\ : InMux
    port map (
            O => \N__4834\,
            I => \N__4826\
        );

    \I__924\ : InMux
    port map (
            O => \N__4833\,
            I => \N__4823\
        );

    \I__923\ : InMux
    port map (
            O => \N__4832\,
            I => \N__4820\
        );

    \I__922\ : LocalMux
    port map (
            O => \N__4829\,
            I => \N__4817\
        );

    \I__921\ : LocalMux
    port map (
            O => \N__4826\,
            I => \pc.program_counterZ0Z_1\
        );

    \I__920\ : LocalMux
    port map (
            O => \N__4823\,
            I => \pc.program_counterZ0Z_1\
        );

    \I__919\ : LocalMux
    port map (
            O => \N__4820\,
            I => \pc.program_counterZ0Z_1\
        );

    \I__918\ : Odrv12
    port map (
            O => \N__4817\,
            I => \pc.program_counterZ0Z_1\
        );

    \I__917\ : ClkMux
    port map (
            O => \N__4808\,
            I => \N__4700\
        );

    \I__916\ : ClkMux
    port map (
            O => \N__4807\,
            I => \N__4700\
        );

    \I__915\ : ClkMux
    port map (
            O => \N__4806\,
            I => \N__4700\
        );

    \I__914\ : ClkMux
    port map (
            O => \N__4805\,
            I => \N__4700\
        );

    \I__913\ : ClkMux
    port map (
            O => \N__4804\,
            I => \N__4700\
        );

    \I__912\ : ClkMux
    port map (
            O => \N__4803\,
            I => \N__4700\
        );

    \I__911\ : ClkMux
    port map (
            O => \N__4802\,
            I => \N__4700\
        );

    \I__910\ : ClkMux
    port map (
            O => \N__4801\,
            I => \N__4700\
        );

    \I__909\ : ClkMux
    port map (
            O => \N__4800\,
            I => \N__4700\
        );

    \I__908\ : ClkMux
    port map (
            O => \N__4799\,
            I => \N__4700\
        );

    \I__907\ : ClkMux
    port map (
            O => \N__4798\,
            I => \N__4700\
        );

    \I__906\ : ClkMux
    port map (
            O => \N__4797\,
            I => \N__4700\
        );

    \I__905\ : ClkMux
    port map (
            O => \N__4796\,
            I => \N__4700\
        );

    \I__904\ : ClkMux
    port map (
            O => \N__4795\,
            I => \N__4700\
        );

    \I__903\ : ClkMux
    port map (
            O => \N__4794\,
            I => \N__4700\
        );

    \I__902\ : ClkMux
    port map (
            O => \N__4793\,
            I => \N__4700\
        );

    \I__901\ : ClkMux
    port map (
            O => \N__4792\,
            I => \N__4700\
        );

    \I__900\ : ClkMux
    port map (
            O => \N__4791\,
            I => \N__4700\
        );

    \I__899\ : ClkMux
    port map (
            O => \N__4790\,
            I => \N__4700\
        );

    \I__898\ : ClkMux
    port map (
            O => \N__4789\,
            I => \N__4700\
        );

    \I__897\ : ClkMux
    port map (
            O => \N__4788\,
            I => \N__4700\
        );

    \I__896\ : ClkMux
    port map (
            O => \N__4787\,
            I => \N__4700\
        );

    \I__895\ : ClkMux
    port map (
            O => \N__4786\,
            I => \N__4700\
        );

    \I__894\ : ClkMux
    port map (
            O => \N__4785\,
            I => \N__4700\
        );

    \I__893\ : ClkMux
    port map (
            O => \N__4784\,
            I => \N__4700\
        );

    \I__892\ : ClkMux
    port map (
            O => \N__4783\,
            I => \N__4700\
        );

    \I__891\ : ClkMux
    port map (
            O => \N__4782\,
            I => \N__4700\
        );

    \I__890\ : ClkMux
    port map (
            O => \N__4781\,
            I => \N__4700\
        );

    \I__889\ : ClkMux
    port map (
            O => \N__4780\,
            I => \N__4700\
        );

    \I__888\ : ClkMux
    port map (
            O => \N__4779\,
            I => \N__4700\
        );

    \I__887\ : ClkMux
    port map (
            O => \N__4778\,
            I => \N__4700\
        );

    \I__886\ : ClkMux
    port map (
            O => \N__4777\,
            I => \N__4700\
        );

    \I__885\ : ClkMux
    port map (
            O => \N__4776\,
            I => \N__4700\
        );

    \I__884\ : ClkMux
    port map (
            O => \N__4775\,
            I => \N__4700\
        );

    \I__883\ : ClkMux
    port map (
            O => \N__4774\,
            I => \N__4700\
        );

    \I__882\ : ClkMux
    port map (
            O => \N__4773\,
            I => \N__4700\
        );

    \I__881\ : GlobalMux
    port map (
            O => \N__4700\,
            I => \N__4697\
        );

    \I__880\ : gio2CtrlBuf
    port map (
            O => \N__4697\,
            I => buf_clk_1_g
        );

    \I__879\ : CascadeMux
    port map (
            O => \N__4694\,
            I => \N__4687\
        );

    \I__878\ : InMux
    port map (
            O => \N__4693\,
            I => \N__4681\
        );

    \I__877\ : InMux
    port map (
            O => \N__4692\,
            I => \N__4681\
        );

    \I__876\ : InMux
    port map (
            O => \N__4691\,
            I => \N__4678\
        );

    \I__875\ : InMux
    port map (
            O => \N__4690\,
            I => \N__4673\
        );

    \I__874\ : InMux
    port map (
            O => \N__4687\,
            I => \N__4673\
        );

    \I__873\ : CascadeMux
    port map (
            O => \N__4686\,
            I => \N__4670\
        );

    \I__872\ : LocalMux
    port map (
            O => \N__4681\,
            I => \N__4663\
        );

    \I__871\ : LocalMux
    port map (
            O => \N__4678\,
            I => \N__4658\
        );

    \I__870\ : LocalMux
    port map (
            O => \N__4673\,
            I => \N__4658\
        );

    \I__869\ : InMux
    port map (
            O => \N__4670\,
            I => \N__4655\
        );

    \I__868\ : InMux
    port map (
            O => \N__4669\,
            I => \N__4651\
        );

    \I__867\ : CascadeMux
    port map (
            O => \N__4668\,
            I => \N__4648\
        );

    \I__866\ : InMux
    port map (
            O => \N__4667\,
            I => \N__4645\
        );

    \I__865\ : CascadeMux
    port map (
            O => \N__4666\,
            I => \N__4641\
        );

    \I__864\ : Span4Mux_h
    port map (
            O => \N__4663\,
            I => \N__4632\
        );

    \I__863\ : Span4Mux_v
    port map (
            O => \N__4658\,
            I => \N__4632\
        );

    \I__862\ : LocalMux
    port map (
            O => \N__4655\,
            I => \N__4632\
        );

    \I__861\ : CascadeMux
    port map (
            O => \N__4654\,
            I => \N__4629\
        );

    \I__860\ : LocalMux
    port map (
            O => \N__4651\,
            I => \N__4626\
        );

    \I__859\ : InMux
    port map (
            O => \N__4648\,
            I => \N__4623\
        );

    \I__858\ : LocalMux
    port map (
            O => \N__4645\,
            I => \N__4620\
        );

    \I__857\ : InMux
    port map (
            O => \N__4644\,
            I => \N__4615\
        );

    \I__856\ : InMux
    port map (
            O => \N__4641\,
            I => \N__4615\
        );

    \I__855\ : InMux
    port map (
            O => \N__4640\,
            I => \N__4610\
        );

    \I__854\ : InMux
    port map (
            O => \N__4639\,
            I => \N__4610\
        );

    \I__853\ : Span4Mux_h
    port map (
            O => \N__4632\,
            I => \N__4607\
        );

    \I__852\ : InMux
    port map (
            O => \N__4629\,
            I => \N__4604\
        );

    \I__851\ : Odrv4
    port map (
            O => \N__4626\,
            I => \seq_T_2\
        );

    \I__850\ : LocalMux
    port map (
            O => \N__4623\,
            I => \seq_T_2\
        );

    \I__849\ : Odrv12
    port map (
            O => \N__4620\,
            I => \seq_T_2\
        );

    \I__848\ : LocalMux
    port map (
            O => \N__4615\,
            I => \seq_T_2\
        );

    \I__847\ : LocalMux
    port map (
            O => \N__4610\,
            I => \seq_T_2\
        );

    \I__846\ : Odrv4
    port map (
            O => \N__4607\,
            I => \seq_T_2\
        );

    \I__845\ : LocalMux
    port map (
            O => \N__4604\,
            I => \seq_T_2\
        );

    \I__844\ : InMux
    port map (
            O => \N__4589\,
            I => \N__4584\
        );

    \I__843\ : InMux
    port map (
            O => \N__4588\,
            I => \N__4581\
        );

    \I__842\ : InMux
    port map (
            O => \N__4587\,
            I => \N__4574\
        );

    \I__841\ : LocalMux
    port map (
            O => \N__4584\,
            I => \N__4571\
        );

    \I__840\ : LocalMux
    port map (
            O => \N__4581\,
            I => \N__4568\
        );

    \I__839\ : InMux
    port map (
            O => \N__4580\,
            I => \N__4563\
        );

    \I__838\ : InMux
    port map (
            O => \N__4579\,
            I => \N__4563\
        );

    \I__837\ : InMux
    port map (
            O => \N__4578\,
            I => \N__4558\
        );

    \I__836\ : InMux
    port map (
            O => \N__4577\,
            I => \N__4558\
        );

    \I__835\ : LocalMux
    port map (
            O => \N__4574\,
            I => \N__4555\
        );

    \I__834\ : Span4Mux_v
    port map (
            O => \N__4571\,
            I => \N__4548\
        );

    \I__833\ : Span4Mux_v
    port map (
            O => \N__4568\,
            I => \N__4548\
        );

    \I__832\ : LocalMux
    port map (
            O => \N__4563\,
            I => \N__4548\
        );

    \I__831\ : LocalMux
    port map (
            O => \N__4558\,
            I => \N__4544\
        );

    \I__830\ : Span4Mux_s2_v
    port map (
            O => \N__4555\,
            I => \N__4536\
        );

    \I__829\ : Span4Mux_h
    port map (
            O => \N__4548\,
            I => \N__4533\
        );

    \I__828\ : InMux
    port map (
            O => \N__4547\,
            I => \N__4530\
        );

    \I__827\ : Span4Mux_h
    port map (
            O => \N__4544\,
            I => \N__4527\
        );

    \I__826\ : InMux
    port map (
            O => \N__4543\,
            I => \N__4522\
        );

    \I__825\ : InMux
    port map (
            O => \N__4542\,
            I => \N__4522\
        );

    \I__824\ : InMux
    port map (
            O => \N__4541\,
            I => \N__4515\
        );

    \I__823\ : InMux
    port map (
            O => \N__4540\,
            I => \N__4515\
        );

    \I__822\ : InMux
    port map (
            O => \N__4539\,
            I => \N__4515\
        );

    \I__821\ : Odrv4
    port map (
            O => \N__4536\,
            I => \seq_PC_LD_0_0\
        );

    \I__820\ : Odrv4
    port map (
            O => \N__4533\,
            I => \seq_PC_LD_0_0\
        );

    \I__819\ : LocalMux
    port map (
            O => \N__4530\,
            I => \seq_PC_LD_0_0\
        );

    \I__818\ : Odrv4
    port map (
            O => \N__4527\,
            I => \seq_PC_LD_0_0\
        );

    \I__817\ : LocalMux
    port map (
            O => \N__4522\,
            I => \seq_PC_LD_0_0\
        );

    \I__816\ : LocalMux
    port map (
            O => \N__4515\,
            I => \seq_PC_LD_0_0\
        );

    \I__815\ : InMux
    port map (
            O => \N__4502\,
            I => \N__4498\
        );

    \I__814\ : InMux
    port map (
            O => \N__4501\,
            I => \N__4494\
        );

    \I__813\ : LocalMux
    port map (
            O => \N__4498\,
            I => \N__4489\
        );

    \I__812\ : InMux
    port map (
            O => \N__4497\,
            I => \N__4486\
        );

    \I__811\ : LocalMux
    port map (
            O => \N__4494\,
            I => \N__4482\
        );

    \I__810\ : InMux
    port map (
            O => \N__4493\,
            I => \N__4479\
        );

    \I__809\ : InMux
    port map (
            O => \N__4492\,
            I => \N__4476\
        );

    \I__808\ : Span4Mux_v
    port map (
            O => \N__4489\,
            I => \N__4473\
        );

    \I__807\ : LocalMux
    port map (
            O => \N__4486\,
            I => \N__4470\
        );

    \I__806\ : InMux
    port map (
            O => \N__4485\,
            I => \N__4467\
        );

    \I__805\ : Span4Mux_v
    port map (
            O => \N__4482\,
            I => \N__4462\
        );

    \I__804\ : LocalMux
    port map (
            O => \N__4479\,
            I => \N__4462\
        );

    \I__803\ : LocalMux
    port map (
            O => \N__4476\,
            I => \N__4459\
        );

    \I__802\ : Span4Mux_v
    port map (
            O => \N__4473\,
            I => \N__4454\
        );

    \I__801\ : Span4Mux_v
    port map (
            O => \N__4470\,
            I => \N__4447\
        );

    \I__800\ : LocalMux
    port map (
            O => \N__4467\,
            I => \N__4447\
        );

    \I__799\ : Span4Mux_h
    port map (
            O => \N__4462\,
            I => \N__4447\
        );

    \I__798\ : Span4Mux_h
    port map (
            O => \N__4459\,
            I => \N__4444\
        );

    \I__797\ : InMux
    port map (
            O => \N__4458\,
            I => \N__4439\
        );

    \I__796\ : InMux
    port map (
            O => \N__4457\,
            I => \N__4439\
        );

    \I__795\ : Odrv4
    port map (
            O => \N__4454\,
            I => \seq_MAR_LD_2\
        );

    \I__794\ : Odrv4
    port map (
            O => \N__4447\,
            I => \seq_MAR_LD_2\
        );

    \I__793\ : Odrv4
    port map (
            O => \N__4444\,
            I => \seq_MAR_LD_2\
        );

    \I__792\ : LocalMux
    port map (
            O => \N__4439\,
            I => \seq_MAR_LD_2\
        );

    \I__791\ : CascadeMux
    port map (
            O => \N__4430\,
            I => \N__4427\
        );

    \I__790\ : InMux
    port map (
            O => \N__4427\,
            I => \N__4424\
        );

    \I__789\ : LocalMux
    port map (
            O => \N__4424\,
            I => \N__4421\
        );

    \I__788\ : Odrv4
    port map (
            O => \N__4421\,
            I => \seq.gZ0Z2\
        );

    \I__787\ : InMux
    port map (
            O => \N__4418\,
            I => \N__4414\
        );

    \I__786\ : InMux
    port map (
            O => \N__4417\,
            I => \N__4408\
        );

    \I__785\ : LocalMux
    port map (
            O => \N__4414\,
            I => \N__4405\
        );

    \I__784\ : InMux
    port map (
            O => \N__4413\,
            I => \N__4402\
        );

    \I__783\ : InMux
    port map (
            O => \N__4412\,
            I => \N__4397\
        );

    \I__782\ : InMux
    port map (
            O => \N__4411\,
            I => \N__4397\
        );

    \I__781\ : LocalMux
    port map (
            O => \N__4408\,
            I => ir_out_5
        );

    \I__780\ : Odrv4
    port map (
            O => \N__4405\,
            I => ir_out_5
        );

    \I__779\ : LocalMux
    port map (
            O => \N__4402\,
            I => ir_out_5
        );

    \I__778\ : LocalMux
    port map (
            O => \N__4397\,
            I => ir_out_5
        );

    \I__777\ : InMux
    port map (
            O => \N__4388\,
            I => \N__4384\
        );

    \I__776\ : InMux
    port map (
            O => \N__4387\,
            I => \N__4380\
        );

    \I__775\ : LocalMux
    port map (
            O => \N__4384\,
            I => \N__4377\
        );

    \I__774\ : InMux
    port map (
            O => \N__4383\,
            I => \N__4374\
        );

    \I__773\ : LocalMux
    port map (
            O => \N__4380\,
            I => \N__4369\
        );

    \I__772\ : Span4Mux_h
    port map (
            O => \N__4377\,
            I => \N__4369\
        );

    \I__771\ : LocalMux
    port map (
            O => \N__4374\,
            I => \N__4366\
        );

    \I__770\ : Span4Mux_v
    port map (
            O => \N__4369\,
            I => \N__4363\
        );

    \I__769\ : Odrv4
    port map (
            O => \N__4366\,
            I => bus_7
        );

    \I__768\ : Odrv4
    port map (
            O => \N__4363\,
            I => bus_7
        );

    \I__767\ : InMux
    port map (
            O => \N__4358\,
            I => \N__4355\
        );

    \I__766\ : LocalMux
    port map (
            O => \N__4355\,
            I => \N__4352\
        );

    \I__765\ : Span4Mux_s2_v
    port map (
            O => \N__4352\,
            I => \N__4348\
        );

    \I__764\ : InMux
    port map (
            O => \N__4351\,
            I => \N__4345\
        );

    \I__763\ : Odrv4
    port map (
            O => \N__4348\,
            I => \N_5_0\
        );

    \I__762\ : LocalMux
    port map (
            O => \N__4345\,
            I => \N_5_0\
        );

    \I__761\ : CascadeMux
    port map (
            O => \N__4340\,
            I => \N_1_0_cascade_\
        );

    \I__760\ : InMux
    port map (
            O => \N__4337\,
            I => \N__4334\
        );

    \I__759\ : LocalMux
    port map (
            O => \N__4334\,
            I => \N__4331\
        );

    \I__758\ : Span4Mux_v
    port map (
            O => \N__4331\,
            I => \N__4328\
        );

    \I__757\ : Span4Mux_v
    port map (
            O => \N__4328\,
            I => \N__4325\
        );

    \I__756\ : Odrv4
    port map (
            O => \N__4325\,
            I => \seq_un1_HLT_0\
        );

    \I__755\ : InMux
    port map (
            O => \N__4322\,
            I => \N__4319\
        );

    \I__754\ : LocalMux
    port map (
            O => \N__4319\,
            I => \seq.un1_HLT_1_reti\
        );

    \I__753\ : InMux
    port map (
            O => \N__4316\,
            I => \N__4313\
        );

    \I__752\ : LocalMux
    port map (
            O => \N__4313\,
            I => \N__4310\
        );

    \I__751\ : Span4Mux_s3_h
    port map (
            O => \N__4310\,
            I => \N__4305\
        );

    \I__750\ : InMux
    port map (
            O => \N__4309\,
            I => \N__4302\
        );

    \I__749\ : InMux
    port map (
            O => \N__4308\,
            I => \N__4299\
        );

    \I__748\ : Odrv4
    port map (
            O => \N__4305\,
            I => \N_2_0\
        );

    \I__747\ : LocalMux
    port map (
            O => \N__4302\,
            I => \N_2_0\
        );

    \I__746\ : LocalMux
    port map (
            O => \N__4299\,
            I => \N_2_0\
        );

    \I__745\ : CascadeMux
    port map (
            O => \N__4292\,
            I => \N__4289\
        );

    \I__744\ : InMux
    port map (
            O => \N__4289\,
            I => \N__4286\
        );

    \I__743\ : LocalMux
    port map (
            O => \N__4286\,
            I => \N__4283\
        );

    \I__742\ : Span4Mux_v
    port map (
            O => \N__4283\,
            I => \N__4280\
        );

    \I__741\ : Odrv4
    port map (
            O => \N__4280\,
            I => \seq.un1_HLT_1\
        );

    \I__740\ : CascadeMux
    port map (
            O => \N__4277\,
            I => \bus_1_cascade_\
        );

    \I__739\ : InMux
    port map (
            O => \N__4274\,
            I => \N__4268\
        );

    \I__738\ : InMux
    port map (
            O => \N__4273\,
            I => \N__4264\
        );

    \I__737\ : InMux
    port map (
            O => \N__4272\,
            I => \N__4259\
        );

    \I__736\ : InMux
    port map (
            O => \N__4271\,
            I => \N__4259\
        );

    \I__735\ : LocalMux
    port map (
            O => \N__4268\,
            I => \N__4256\
        );

    \I__734\ : InMux
    port map (
            O => \N__4267\,
            I => \N__4253\
        );

    \I__733\ : LocalMux
    port map (
            O => \N__4264\,
            I => \N__4243\
        );

    \I__732\ : LocalMux
    port map (
            O => \N__4259\,
            I => \N__4243\
        );

    \I__731\ : Span4Mux_v
    port map (
            O => \N__4256\,
            I => \N__4238\
        );

    \I__730\ : LocalMux
    port map (
            O => \N__4253\,
            I => \N__4238\
        );

    \I__729\ : InMux
    port map (
            O => \N__4252\,
            I => \N__4233\
        );

    \I__728\ : InMux
    port map (
            O => \N__4251\,
            I => \N__4233\
        );

    \I__727\ : InMux
    port map (
            O => \N__4250\,
            I => \N__4228\
        );

    \I__726\ : InMux
    port map (
            O => \N__4249\,
            I => \N__4228\
        );

    \I__725\ : InMux
    port map (
            O => \N__4248\,
            I => \N__4225\
        );

    \I__724\ : Odrv4
    port map (
            O => \N__4243\,
            I => \seq_D_6\
        );

    \I__723\ : Odrv4
    port map (
            O => \N__4238\,
            I => \seq_D_6\
        );

    \I__722\ : LocalMux
    port map (
            O => \N__4233\,
            I => \seq_D_6\
        );

    \I__721\ : LocalMux
    port map (
            O => \N__4228\,
            I => \seq_D_6\
        );

    \I__720\ : LocalMux
    port map (
            O => \N__4225\,
            I => \seq_D_6\
        );

    \I__719\ : InMux
    port map (
            O => \N__4214\,
            I => \N__4210\
        );

    \I__718\ : InMux
    port map (
            O => \N__4213\,
            I => \N__4207\
        );

    \I__717\ : LocalMux
    port map (
            O => \N__4210\,
            I => \N__4198\
        );

    \I__716\ : LocalMux
    port map (
            O => \N__4207\,
            I => \N__4198\
        );

    \I__715\ : InMux
    port map (
            O => \N__4206\,
            I => \N__4195\
        );

    \I__714\ : InMux
    port map (
            O => \N__4205\,
            I => \N__4191\
        );

    \I__713\ : InMux
    port map (
            O => \N__4204\,
            I => \N__4188\
        );

    \I__712\ : InMux
    port map (
            O => \N__4203\,
            I => \N__4185\
        );

    \I__711\ : Span4Mux_h
    port map (
            O => \N__4198\,
            I => \N__4180\
        );

    \I__710\ : LocalMux
    port map (
            O => \N__4195\,
            I => \N__4176\
        );

    \I__709\ : InMux
    port map (
            O => \N__4194\,
            I => \N__4173\
        );

    \I__708\ : LocalMux
    port map (
            O => \N__4191\,
            I => \N__4166\
        );

    \I__707\ : LocalMux
    port map (
            O => \N__4188\,
            I => \N__4166\
        );

    \I__706\ : LocalMux
    port map (
            O => \N__4185\,
            I => \N__4166\
        );

    \I__705\ : InMux
    port map (
            O => \N__4184\,
            I => \N__4161\
        );

    \I__704\ : InMux
    port map (
            O => \N__4183\,
            I => \N__4161\
        );

    \I__703\ : Span4Mux_v
    port map (
            O => \N__4180\,
            I => \N__4158\
        );

    \I__702\ : InMux
    port map (
            O => \N__4179\,
            I => \N__4155\
        );

    \I__701\ : Span4Mux_h
    port map (
            O => \N__4176\,
            I => \N__4150\
        );

    \I__700\ : LocalMux
    port map (
            O => \N__4173\,
            I => \N__4150\
        );

    \I__699\ : Span4Mux_v
    port map (
            O => \N__4166\,
            I => \N__4147\
        );

    \I__698\ : LocalMux
    port map (
            O => \N__4161\,
            I => \T_0_fast_RNILB791_2\
        );

    \I__697\ : Odrv4
    port map (
            O => \N__4158\,
            I => \T_0_fast_RNILB791_2\
        );

    \I__696\ : LocalMux
    port map (
            O => \N__4155\,
            I => \T_0_fast_RNILB791_2\
        );

    \I__695\ : Odrv4
    port map (
            O => \N__4150\,
            I => \T_0_fast_RNILB791_2\
        );

    \I__694\ : Odrv4
    port map (
            O => \N__4147\,
            I => \T_0_fast_RNILB791_2\
        );

    \I__693\ : CascadeMux
    port map (
            O => \N__4136\,
            I => \N__4132\
        );

    \I__692\ : InMux
    port map (
            O => \N__4135\,
            I => \N__4129\
        );

    \I__691\ : InMux
    port map (
            O => \N__4132\,
            I => \N__4126\
        );

    \I__690\ : LocalMux
    port map (
            O => \N__4129\,
            I => \AR_out_1\
        );

    \I__689\ : LocalMux
    port map (
            O => \N__4126\,
            I => \AR_out_1\
        );

    \I__688\ : CascadeMux
    port map (
            O => \N__4121\,
            I => \ALU_main_N_44_0_cascade_\
        );

    \I__687\ : InMux
    port map (
            O => \N__4118\,
            I => \N__4112\
        );

    \I__686\ : InMux
    port map (
            O => \N__4117\,
            I => \N__4112\
        );

    \I__685\ : LocalMux
    port map (
            O => \N__4112\,
            I => \un1_A_cry_2_c_RNI1TTO2\
        );

    \I__684\ : InMux
    port map (
            O => \N__4109\,
            I => \N__4106\
        );

    \I__683\ : LocalMux
    port map (
            O => \N__4106\,
            I => \N__4103\
        );

    \I__682\ : Odrv4
    port map (
            O => \N__4103\,
            I => \pc.N_10_i\
        );

    \I__681\ : InMux
    port map (
            O => \N__4100\,
            I => \N__4097\
        );

    \I__680\ : LocalMux
    port map (
            O => \N__4097\,
            I => \N__4094\
        );

    \I__679\ : Span12Mux_s4_v
    port map (
            O => \N__4094\,
            I => \N__4091\
        );

    \I__678\ : Odrv12
    port map (
            O => \N__4091\,
            I => \pc.G_10_0_1_1\
        );

    \I__677\ : InMux
    port map (
            O => \N__4088\,
            I => \N__4085\
        );

    \I__676\ : LocalMux
    port map (
            O => \N__4085\,
            I => \N__4082\
        );

    \I__675\ : Odrv4
    port map (
            O => \N__4082\,
            I => \pc.G_10_0_1\
        );

    \I__674\ : CascadeMux
    port map (
            O => \N__4079\,
            I => \N__4076\
        );

    \I__673\ : InMux
    port map (
            O => \N__4076\,
            I => \N__4073\
        );

    \I__672\ : LocalMux
    port map (
            O => \N__4073\,
            I => \ALU_main_N_44_1\
        );

    \I__671\ : InMux
    port map (
            O => \N__4070\,
            I => \N__4067\
        );

    \I__670\ : LocalMux
    port map (
            O => \N__4067\,
            I => \N__4064\
        );

    \I__669\ : Odrv12
    port map (
            O => \N__4064\,
            I => \pc.un1_inc_0_0\
        );

    \I__668\ : InMux
    port map (
            O => \N__4061\,
            I => \N__4058\
        );

    \I__667\ : LocalMux
    port map (
            O => \N__4058\,
            I => \N__4055\
        );

    \I__666\ : Span4Mux_v
    port map (
            O => \N__4055\,
            I => \N__4052\
        );

    \I__665\ : Odrv4
    port map (
            O => \N__4052\,
            I => \pc.out_1_iv_1_1\
        );

    \I__664\ : CascadeMux
    port map (
            O => \N__4049\,
            I => \N__4046\
        );

    \I__663\ : InMux
    port map (
            O => \N__4046\,
            I => \N__4043\
        );

    \I__662\ : LocalMux
    port map (
            O => \N__4043\,
            I => \N__4040\
        );

    \I__661\ : Span4Mux_v
    port map (
            O => \N__4040\,
            I => \N__4037\
        );

    \I__660\ : Span4Mux_h
    port map (
            O => \N__4037\,
            I => \N__4034\
        );

    \I__659\ : Odrv4
    port map (
            O => \N__4034\,
            I => \mem_data_2_7_0__N_16_0\
        );

    \I__658\ : InMux
    port map (
            O => \N__4031\,
            I => \N__4028\
        );

    \I__657\ : LocalMux
    port map (
            O => \N__4028\,
            I => \N__4025\
        );

    \I__656\ : Span4Mux_h
    port map (
            O => \N__4025\,
            I => \N__4022\
        );

    \I__655\ : Odrv4
    port map (
            O => \N__4022\,
            I => \pc.g0_rn_1\
        );

    \I__654\ : CascadeMux
    port map (
            O => \N__4019\,
            I => \pc.g0_sn_cascade_\
        );

    \I__653\ : InMux
    port map (
            O => \N__4016\,
            I => \N__4013\
        );

    \I__652\ : LocalMux
    port map (
            O => \N__4013\,
            I => alu_out_m_0_3
        );

    \I__651\ : InMux
    port map (
            O => \N__4010\,
            I => \N__4006\
        );

    \I__650\ : InMux
    port map (
            O => \N__4009\,
            I => \N__4003\
        );

    \I__649\ : LocalMux
    port map (
            O => \N__4006\,
            I => \N__4000\
        );

    \I__648\ : LocalMux
    port map (
            O => \N__4003\,
            I => \N__3997\
        );

    \I__647\ : Span4Mux_v
    port map (
            O => \N__4000\,
            I => \N__3992\
        );

    \I__646\ : Span4Mux_s3_h
    port map (
            O => \N__3997\,
            I => \N__3992\
        );

    \I__645\ : Odrv4
    port map (
            O => \N__3992\,
            I => \pc.program_counterZ0Z_3\
        );

    \I__644\ : InMux
    port map (
            O => \N__3989\,
            I => \N__3986\
        );

    \I__643\ : LocalMux
    port map (
            O => \N__3986\,
            I => \N__3982\
        );

    \I__642\ : InMux
    port map (
            O => \N__3985\,
            I => \N__3979\
        );

    \I__641\ : Span4Mux_h
    port map (
            O => \N__3982\,
            I => \N__3976\
        );

    \I__640\ : LocalMux
    port map (
            O => \N__3979\,
            I => \seq_un1_AR_OE_0_0\
        );

    \I__639\ : Odrv4
    port map (
            O => \N__3976\,
            I => \seq_un1_AR_OE_0_0\
        );

    \I__638\ : InMux
    port map (
            O => \N__3971\,
            I => \N__3968\
        );

    \I__637\ : LocalMux
    port map (
            O => \N__3968\,
            I => \N__3960\
        );

    \I__636\ : InMux
    port map (
            O => \N__3967\,
            I => \N__3955\
        );

    \I__635\ : InMux
    port map (
            O => \N__3966\,
            I => \N__3955\
        );

    \I__634\ : CascadeMux
    port map (
            O => \N__3965\,
            I => \N__3952\
        );

    \I__633\ : InMux
    port map (
            O => \N__3964\,
            I => \N__3949\
        );

    \I__632\ : InMux
    port map (
            O => \N__3963\,
            I => \N__3946\
        );

    \I__631\ : Span4Mux_v
    port map (
            O => \N__3960\,
            I => \N__3943\
        );

    \I__630\ : LocalMux
    port map (
            O => \N__3955\,
            I => \N__3940\
        );

    \I__629\ : InMux
    port map (
            O => \N__3952\,
            I => \N__3937\
        );

    \I__628\ : LocalMux
    port map (
            O => \N__3949\,
            I => ir_out_6
        );

    \I__627\ : LocalMux
    port map (
            O => \N__3946\,
            I => ir_out_6
        );

    \I__626\ : Odrv4
    port map (
            O => \N__3943\,
            I => ir_out_6
        );

    \I__625\ : Odrv12
    port map (
            O => \N__3940\,
            I => ir_out_6
        );

    \I__624\ : LocalMux
    port map (
            O => \N__3937\,
            I => ir_out_6
        );

    \I__623\ : InMux
    port map (
            O => \N__3926\,
            I => \N__3922\
        );

    \I__622\ : CascadeMux
    port map (
            O => \N__3925\,
            I => \N__3919\
        );

    \I__621\ : LocalMux
    port map (
            O => \N__3922\,
            I => \N__3916\
        );

    \I__620\ : InMux
    port map (
            O => \N__3919\,
            I => \N__3913\
        );

    \I__619\ : Span4Mux_s1_v
    port map (
            O => \N__3916\,
            I => \N__3909\
        );

    \I__618\ : LocalMux
    port map (
            O => \N__3913\,
            I => \N__3906\
        );

    \I__617\ : InMux
    port map (
            O => \N__3912\,
            I => \N__3903\
        );

    \I__616\ : Span4Mux_v
    port map (
            O => \N__3909\,
            I => \N__3900\
        );

    \I__615\ : Span4Mux_h
    port map (
            O => \N__3906\,
            I => \N__3897\
        );

    \I__614\ : LocalMux
    port map (
            O => \N__3903\,
            I => \AR.ff4.AR_out_3\
        );

    \I__613\ : Odrv4
    port map (
            O => \N__3900\,
            I => \AR.ff4.AR_out_3\
        );

    \I__612\ : Odrv4
    port map (
            O => \N__3897\,
            I => \AR.ff4.AR_out_3\
        );

    \I__611\ : InMux
    port map (
            O => \N__3890\,
            I => \N__3885\
        );

    \I__610\ : InMux
    port map (
            O => \N__3889\,
            I => \N__3882\
        );

    \I__609\ : InMux
    port map (
            O => \N__3888\,
            I => \N__3879\
        );

    \I__608\ : LocalMux
    port map (
            O => \N__3885\,
            I => \N__3876\
        );

    \I__607\ : LocalMux
    port map (
            O => \N__3882\,
            I => \N__3872\
        );

    \I__606\ : LocalMux
    port map (
            O => \N__3879\,
            I => \N__3869\
        );

    \I__605\ : Span4Mux_v
    port map (
            O => \N__3876\,
            I => \N__3866\
        );

    \I__604\ : InMux
    port map (
            O => \N__3875\,
            I => \N__3863\
        );

    \I__603\ : Span4Mux_h
    port map (
            O => \N__3872\,
            I => \N__3860\
        );

    \I__602\ : Span4Mux_s2_h
    port map (
            O => \N__3869\,
            I => \N__3857\
        );

    \I__601\ : Odrv4
    port map (
            O => \N__3866\,
            I => ir_out_3
        );

    \I__600\ : LocalMux
    port map (
            O => \N__3863\,
            I => ir_out_3
        );

    \I__599\ : Odrv4
    port map (
            O => \N__3860\,
            I => ir_out_3
        );

    \I__598\ : Odrv4
    port map (
            O => \N__3857\,
            I => ir_out_3
        );

    \I__597\ : InMux
    port map (
            O => \N__3848\,
            I => \N__3845\
        );

    \I__596\ : LocalMux
    port map (
            O => \N__3845\,
            I => \pc.tbuf.g0_0_1_0\
        );

    \I__595\ : CascadeMux
    port map (
            O => \N__3842\,
            I => \AR_out_m_3_cascade_\
        );

    \I__594\ : InMux
    port map (
            O => \N__3839\,
            I => \N__3836\
        );

    \I__593\ : LocalMux
    port map (
            O => \N__3836\,
            I => \pc.g0_0\
        );

    \I__592\ : CascadeMux
    port map (
            O => \N__3833\,
            I => \N__3830\
        );

    \I__591\ : InMux
    port map (
            O => \N__3830\,
            I => \N__3827\
        );

    \I__590\ : LocalMux
    port map (
            O => \N__3827\,
            I => \ALU_main.un1_A_axb_2_l_ofxZ0\
        );

    \I__589\ : InMux
    port map (
            O => \N__3824\,
            I => \N__3821\
        );

    \I__588\ : LocalMux
    port map (
            O => \N__3821\,
            I => \N__3817\
        );

    \I__587\ : InMux
    port map (
            O => \N__3820\,
            I => \N__3814\
        );

    \I__586\ : Odrv4
    port map (
            O => \N__3817\,
            I => \un1_A_cry_1_c_RNITKPO2\
        );

    \I__585\ : LocalMux
    port map (
            O => \N__3814\,
            I => \un1_A_cry_1_c_RNITKPO2\
        );

    \I__584\ : InMux
    port map (
            O => \N__3809\,
            I => \ALU_main.un1_A_cry_1\
        );

    \I__583\ : InMux
    port map (
            O => \N__3806\,
            I => \ALU_main.un1_A_cry_2\
        );

    \I__582\ : InMux
    port map (
            O => \N__3803\,
            I => \ALU_main.un1_A_cry_3\
        );

    \I__581\ : InMux
    port map (
            O => \N__3800\,
            I => \ALU_main.un1_A_cry_4\
        );

    \I__580\ : InMux
    port map (
            O => \N__3797\,
            I => \ALU_main.un1_A_cry_5\
        );

    \I__579\ : InMux
    port map (
            O => \N__3794\,
            I => \bfn_4_13_0_\
        );

    \I__578\ : InMux
    port map (
            O => \N__3791\,
            I => \N__3788\
        );

    \I__577\ : LocalMux
    port map (
            O => \N__3788\,
            I => \N__3785\
        );

    \I__576\ : Span4Mux_s3_h
    port map (
            O => \N__3785\,
            I => \N__3782\
        );

    \I__575\ : Odrv4
    port map (
            O => \N__3782\,
            I => \ALU_main.un1_A_cry_6_c_RNIP89EZ0Z2\
        );

    \I__574\ : InMux
    port map (
            O => \N__3779\,
            I => \N__3776\
        );

    \I__573\ : LocalMux
    port map (
            O => \N__3776\,
            I => \ALU_main.un1_A_cry_5_c_RNIDLAPZ0Z2\
        );

    \I__572\ : InMux
    port map (
            O => \N__3773\,
            I => \N__3770\
        );

    \I__571\ : LocalMux
    port map (
            O => \N__3770\,
            I => \N__3766\
        );

    \I__570\ : InMux
    port map (
            O => \N__3769\,
            I => \N__3763\
        );

    \I__569\ : Span4Mux_h
    port map (
            O => \N__3766\,
            I => \N__3760\
        );

    \I__568\ : LocalMux
    port map (
            O => \N__3763\,
            I => \N__3757\
        );

    \I__567\ : Odrv4
    port map (
            O => \N__3760\,
            I => \N_30\
        );

    \I__566\ : Odrv4
    port map (
            O => \N__3757\,
            I => \N_30\
        );

    \I__565\ : CascadeMux
    port map (
            O => \N__3752\,
            I => \pc.G_10_0_1_0_cascade_\
        );

    \I__564\ : InMux
    port map (
            O => \N__3749\,
            I => \N__3746\
        );

    \I__563\ : LocalMux
    port map (
            O => \N__3746\,
            I => \N__3743\
        );

    \I__562\ : Odrv4
    port map (
            O => \N__3743\,
            I => \pc.G_10_0_sx\
        );

    \I__561\ : CascadeMux
    port map (
            O => \N__3740\,
            I => \N__3737\
        );

    \I__560\ : InMux
    port map (
            O => \N__3737\,
            I => \N__3734\
        );

    \I__559\ : LocalMux
    port map (
            O => \N__3734\,
            I => \pc.G_10_0_5_1\
        );

    \I__558\ : InMux
    port map (
            O => \N__3731\,
            I => \N__3728\
        );

    \I__557\ : LocalMux
    port map (
            O => \N__3728\,
            I => \N__3725\
        );

    \I__556\ : Odrv4
    port map (
            O => \N__3725\,
            I => \ALU_main_N_43_0\
        );

    \I__555\ : CascadeMux
    port map (
            O => \N__3722\,
            I => \N__3719\
        );

    \I__554\ : InMux
    port map (
            O => \N__3719\,
            I => \N__3715\
        );

    \I__553\ : InMux
    port map (
            O => \N__3718\,
            I => \N__3712\
        );

    \I__552\ : LocalMux
    port map (
            O => \N__3715\,
            I => \N__3708\
        );

    \I__551\ : LocalMux
    port map (
            O => \N__3712\,
            I => \N__3705\
        );

    \I__550\ : InMux
    port map (
            O => \N__3711\,
            I => \N__3701\
        );

    \I__549\ : Span4Mux_v
    port map (
            O => \N__3708\,
            I => \N__3695\
        );

    \I__548\ : Span4Mux_v
    port map (
            O => \N__3705\,
            I => \N__3695\
        );

    \I__547\ : InMux
    port map (
            O => \N__3704\,
            I => \N__3692\
        );

    \I__546\ : LocalMux
    port map (
            O => \N__3701\,
            I => \N__3689\
        );

    \I__545\ : InMux
    port map (
            O => \N__3700\,
            I => \N__3686\
        );

    \I__544\ : Span4Mux_h
    port map (
            O => \N__3695\,
            I => \N__3681\
        );

    \I__543\ : LocalMux
    port map (
            O => \N__3692\,
            I => \N__3681\
        );

    \I__542\ : Span4Mux_s3_h
    port map (
            O => \N__3689\,
            I => \N__3678\
        );

    \I__541\ : LocalMux
    port map (
            O => \N__3686\,
            I => \pc.program_counterZ0Z_2\
        );

    \I__540\ : Odrv4
    port map (
            O => \N__3681\,
            I => \pc.program_counterZ0Z_2\
        );

    \I__539\ : Odrv4
    port map (
            O => \N__3678\,
            I => \pc.program_counterZ0Z_2\
        );

    \I__538\ : InMux
    port map (
            O => \N__3671\,
            I => \N__3667\
        );

    \I__537\ : InMux
    port map (
            O => \N__3670\,
            I => \N__3663\
        );

    \I__536\ : LocalMux
    port map (
            O => \N__3667\,
            I => \N__3659\
        );

    \I__535\ : InMux
    port map (
            O => \N__3666\,
            I => \N__3656\
        );

    \I__534\ : LocalMux
    port map (
            O => \N__3663\,
            I => \N__3653\
        );

    \I__533\ : InMux
    port map (
            O => \N__3662\,
            I => \N__3650\
        );

    \I__532\ : Span4Mux_h
    port map (
            O => \N__3659\,
            I => \N__3645\
        );

    \I__531\ : LocalMux
    port map (
            O => \N__3656\,
            I => \N__3645\
        );

    \I__530\ : Span4Mux_v
    port map (
            O => \N__3653\,
            I => \N__3636\
        );

    \I__529\ : LocalMux
    port map (
            O => \N__3650\,
            I => \N__3636\
        );

    \I__528\ : Span4Mux_v
    port map (
            O => \N__3645\,
            I => \N__3636\
        );

    \I__527\ : InMux
    port map (
            O => \N__3644\,
            I => \N__3631\
        );

    \I__526\ : InMux
    port map (
            O => \N__3643\,
            I => \N__3631\
        );

    \I__525\ : Odrv4
    port map (
            O => \N__3636\,
            I => \pc.program_counterZ0Z_0\
        );

    \I__524\ : LocalMux
    port map (
            O => \N__3631\,
            I => \pc.program_counterZ0Z_0\
        );

    \I__523\ : CascadeMux
    port map (
            O => \N__3626\,
            I => \N__3623\
        );

    \I__522\ : InMux
    port map (
            O => \N__3623\,
            I => \N__3619\
        );

    \I__521\ : InMux
    port map (
            O => \N__3622\,
            I => \N__3616\
        );

    \I__520\ : LocalMux
    port map (
            O => \N__3619\,
            I => \N__3611\
        );

    \I__519\ : LocalMux
    port map (
            O => \N__3616\,
            I => \N__3611\
        );

    \I__518\ : Odrv4
    port map (
            O => \N__3611\,
            I => \seq_S0_0_i\
        );

    \I__517\ : InMux
    port map (
            O => \N__3608\,
            I => \ALU_main.un1_A_cry_0_c_THRU_CO\
        );

    \I__516\ : InMux
    port map (
            O => \N__3605\,
            I => \ALU_main.un1_A_cry_0\
        );

    \I__515\ : CascadeMux
    port map (
            O => \N__3602\,
            I => \IR_OE_1_cascade_\
        );

    \I__514\ : InMux
    port map (
            O => \N__3599\,
            I => \N__3593\
        );

    \I__513\ : InMux
    port map (
            O => \N__3598\,
            I => \N__3593\
        );

    \I__512\ : LocalMux
    port map (
            O => \N__3593\,
            I => \pc.un1_inc_0\
        );

    \I__511\ : CascadeMux
    port map (
            O => \N__3590\,
            I => \N__3587\
        );

    \I__510\ : InMux
    port map (
            O => \N__3587\,
            I => \N__3584\
        );

    \I__509\ : LocalMux
    port map (
            O => \N__3584\,
            I => \N__3581\
        );

    \I__508\ : Odrv12
    port map (
            O => \N__3581\,
            I => \pc.G_12_i_a3_2_3\
        );

    \I__507\ : InMux
    port map (
            O => \N__3578\,
            I => \N__3575\
        );

    \I__506\ : LocalMux
    port map (
            O => \N__3575\,
            I => \pc.G_12_i_a3_2_1\
        );

    \I__505\ : CascadeMux
    port map (
            O => \N__3572\,
            I => \seq.counter.T8_1_cascade_\
        );

    \I__504\ : CascadeMux
    port map (
            O => \N__3569\,
            I => \N__3566\
        );

    \I__503\ : InMux
    port map (
            O => \N__3566\,
            I => \N__3563\
        );

    \I__502\ : LocalMux
    port map (
            O => \N__3563\,
            I => \pc.g1_0\
        );

    \I__501\ : InMux
    port map (
            O => \N__3560\,
            I => \N__3557\
        );

    \I__500\ : LocalMux
    port map (
            O => \N__3557\,
            I => \N__3554\
        );

    \I__499\ : Span4Mux_s3_h
    port map (
            O => \N__3554\,
            I => \N__3551\
        );

    \I__498\ : Odrv4
    port map (
            O => \N__3551\,
            I => \pc.N_188_0\
        );

    \I__497\ : CascadeMux
    port map (
            O => \N__3548\,
            I => \N__3542\
        );

    \I__496\ : CascadeMux
    port map (
            O => \N__3547\,
            I => \N__3538\
        );

    \I__495\ : InMux
    port map (
            O => \N__3546\,
            I => \N__3534\
        );

    \I__494\ : InMux
    port map (
            O => \N__3545\,
            I => \N__3527\
        );

    \I__493\ : InMux
    port map (
            O => \N__3542\,
            I => \N__3527\
        );

    \I__492\ : InMux
    port map (
            O => \N__3541\,
            I => \N__3527\
        );

    \I__491\ : InMux
    port map (
            O => \N__3538\,
            I => \N__3524\
        );

    \I__490\ : CascadeMux
    port map (
            O => \N__3537\,
            I => \N__3520\
        );

    \I__489\ : LocalMux
    port map (
            O => \N__3534\,
            I => \N__3517\
        );

    \I__488\ : LocalMux
    port map (
            O => \N__3527\,
            I => \N__3511\
        );

    \I__487\ : LocalMux
    port map (
            O => \N__3524\,
            I => \N__3508\
        );

    \I__486\ : InMux
    port map (
            O => \N__3523\,
            I => \N__3503\
        );

    \I__485\ : InMux
    port map (
            O => \N__3520\,
            I => \N__3503\
        );

    \I__484\ : Span4Mux_v
    port map (
            O => \N__3517\,
            I => \N__3500\
        );

    \I__483\ : InMux
    port map (
            O => \N__3516\,
            I => \N__3493\
        );

    \I__482\ : InMux
    port map (
            O => \N__3515\,
            I => \N__3493\
        );

    \I__481\ : InMux
    port map (
            O => \N__3514\,
            I => \N__3493\
        );

    \I__480\ : Span4Mux_v
    port map (
            O => \N__3511\,
            I => \N__3486\
        );

    \I__479\ : Span4Mux_v
    port map (
            O => \N__3508\,
            I => \N__3486\
        );

    \I__478\ : LocalMux
    port map (
            O => \N__3503\,
            I => \N__3486\
        );

    \I__477\ : Odrv4
    port map (
            O => \N__3500\,
            I => \seq_T_0\
        );

    \I__476\ : LocalMux
    port map (
            O => \N__3493\,
            I => \seq_T_0\
        );

    \I__475\ : Odrv4
    port map (
            O => \N__3486\,
            I => \seq_T_0\
        );

    \I__474\ : CascadeMux
    port map (
            O => \N__3479\,
            I => \g0_0_1_cascade_\
        );

    \I__473\ : InMux
    port map (
            O => \N__3476\,
            I => \N__3473\
        );

    \I__472\ : LocalMux
    port map (
            O => \N__3473\,
            I => \N__3470\
        );

    \I__471\ : Odrv12
    port map (
            O => \N__3470\,
            I => \seq.counter.un7_ACC_LD_0\
        );

    \I__470\ : InMux
    port map (
            O => \N__3467\,
            I => \N__3464\
        );

    \I__469\ : LocalMux
    port map (
            O => \N__3464\,
            I => \seq.un1_ALU_en_0Z0Z_1\
        );

    \I__468\ : CascadeMux
    port map (
            O => \N__3461\,
            I => \seq.counter.un7_ACC_LD_0_cascade_\
        );

    \I__467\ : CascadeMux
    port map (
            O => \N__3458\,
            I => \IR_OE_2_cascade_\
        );

    \I__466\ : InMux
    port map (
            O => \N__3455\,
            I => \N__3452\
        );

    \I__465\ : LocalMux
    port map (
            O => \N__3452\,
            I => \N__3449\
        );

    \I__464\ : Odrv4
    port map (
            O => \N__3449\,
            I => bus_2
        );

    \I__463\ : InMux
    port map (
            O => \N__3446\,
            I => \N__3443\
        );

    \I__462\ : LocalMux
    port map (
            O => \N__3443\,
            I => \N__3440\
        );

    \I__461\ : Span4Mux_h
    port map (
            O => \N__3440\,
            I => \N__3437\
        );

    \I__460\ : Odrv4
    port map (
            O => \N__3437\,
            I => \seq.g2Z0Z_0\
        );

    \I__459\ : InMux
    port map (
            O => \N__3434\,
            I => \N__3429\
        );

    \I__458\ : CascadeMux
    port map (
            O => \N__3433\,
            I => \N__3425\
        );

    \I__457\ : CascadeMux
    port map (
            O => \N__3432\,
            I => \N__3421\
        );

    \I__456\ : LocalMux
    port map (
            O => \N__3429\,
            I => \N__3418\
        );

    \I__455\ : InMux
    port map (
            O => \N__3428\,
            I => \N__3413\
        );

    \I__454\ : InMux
    port map (
            O => \N__3425\,
            I => \N__3413\
        );

    \I__453\ : CascadeMux
    port map (
            O => \N__3424\,
            I => \N__3410\
        );

    \I__452\ : InMux
    port map (
            O => \N__3421\,
            I => \N__3406\
        );

    \I__451\ : Span4Mux_s1_h
    port map (
            O => \N__3418\,
            I => \N__3401\
        );

    \I__450\ : LocalMux
    port map (
            O => \N__3413\,
            I => \N__3401\
        );

    \I__449\ : InMux
    port map (
            O => \N__3410\,
            I => \N__3398\
        );

    \I__448\ : InMux
    port map (
            O => \N__3409\,
            I => \N__3395\
        );

    \I__447\ : LocalMux
    port map (
            O => \N__3406\,
            I => ir_out_fast_7
        );

    \I__446\ : Odrv4
    port map (
            O => \N__3401\,
            I => ir_out_fast_7
        );

    \I__445\ : LocalMux
    port map (
            O => \N__3398\,
            I => ir_out_fast_7
        );

    \I__444\ : LocalMux
    port map (
            O => \N__3395\,
            I => ir_out_fast_7
        );

    \I__443\ : InMux
    port map (
            O => \N__3386\,
            I => \N__3383\
        );

    \I__442\ : LocalMux
    port map (
            O => \N__3383\,
            I => \N__3380\
        );

    \I__441\ : Odrv4
    port map (
            O => \N__3380\,
            I => \seq.S0_0_i_N_3LZ0Z3\
        );

    \I__440\ : InMux
    port map (
            O => \N__3377\,
            I => \N__3371\
        );

    \I__439\ : InMux
    port map (
            O => \N__3376\,
            I => \N__3366\
        );

    \I__438\ : InMux
    port map (
            O => \N__3375\,
            I => \N__3366\
        );

    \I__437\ : InMux
    port map (
            O => \N__3374\,
            I => \N__3363\
        );

    \I__436\ : LocalMux
    port map (
            O => \N__3371\,
            I => ir_out_i_2_6
        );

    \I__435\ : LocalMux
    port map (
            O => \N__3366\,
            I => ir_out_i_2_6
        );

    \I__434\ : LocalMux
    port map (
            O => \N__3363\,
            I => ir_out_i_2_6
        );

    \I__433\ : InMux
    port map (
            O => \N__3356\,
            I => \N__3352\
        );

    \I__432\ : CascadeMux
    port map (
            O => \N__3355\,
            I => \N__3348\
        );

    \I__431\ : LocalMux
    port map (
            O => \N__3352\,
            I => \N__3345\
        );

    \I__430\ : InMux
    port map (
            O => \N__3351\,
            I => \N__3340\
        );

    \I__429\ : InMux
    port map (
            O => \N__3348\,
            I => \N__3340\
        );

    \I__428\ : Odrv4
    port map (
            O => \N__3345\,
            I => \seq.counter.T_fast_2\
        );

    \I__427\ : LocalMux
    port map (
            O => \N__3340\,
            I => \seq.counter.T_fast_2\
        );

    \I__426\ : InMux
    port map (
            O => \N__3335\,
            I => \N__3332\
        );

    \I__425\ : LocalMux
    port map (
            O => \N__3332\,
            I => \N__3329\
        );

    \I__424\ : Span4Mux_v
    port map (
            O => \N__3329\,
            I => \N__3324\
        );

    \I__423\ : InMux
    port map (
            O => \N__3328\,
            I => \N__3319\
        );

    \I__422\ : InMux
    port map (
            O => \N__3327\,
            I => \N__3319\
        );

    \I__421\ : Odrv4
    port map (
            O => \N__3324\,
            I => \seq_un1_IR_OE_4_1\
        );

    \I__420\ : LocalMux
    port map (
            O => \N__3319\,
            I => \seq_un1_IR_OE_4_1\
        );

    \I__419\ : CascadeMux
    port map (
            O => \N__3314\,
            I => \seq.B_LD_0_2_tz_cascade_\
        );

    \I__418\ : InMux
    port map (
            O => \N__3311\,
            I => \N__3308\
        );

    \I__417\ : LocalMux
    port map (
            O => \N__3308\,
            I => \N__3305\
        );

    \I__416\ : Odrv4
    port map (
            O => \N__3305\,
            I => \seq.counter.T_RNIR83I4_0Z0Z_3\
        );

    \I__415\ : InMux
    port map (
            O => \N__3302\,
            I => \N__3298\
        );

    \I__414\ : InMux
    port map (
            O => \N__3301\,
            I => \N__3292\
        );

    \I__413\ : LocalMux
    port map (
            O => \N__3298\,
            I => \N__3289\
        );

    \I__412\ : InMux
    port map (
            O => \N__3297\,
            I => \N__3286\
        );

    \I__411\ : InMux
    port map (
            O => \N__3296\,
            I => \N__3281\
        );

    \I__410\ : InMux
    port map (
            O => \N__3295\,
            I => \N__3281\
        );

    \I__409\ : LocalMux
    port map (
            O => \N__3292\,
            I => \IR_ff6_q_0_fast\
        );

    \I__408\ : Odrv12
    port map (
            O => \N__3289\,
            I => \IR_ff6_q_0_fast\
        );

    \I__407\ : LocalMux
    port map (
            O => \N__3286\,
            I => \IR_ff6_q_0_fast\
        );

    \I__406\ : LocalMux
    port map (
            O => \N__3281\,
            I => \IR_ff6_q_0_fast\
        );

    \I__405\ : InMux
    port map (
            O => \N__3272\,
            I => \N__3269\
        );

    \I__404\ : LocalMux
    port map (
            O => \N__3269\,
            I => \N__3262\
        );

    \I__403\ : InMux
    port map (
            O => \N__3268\,
            I => \N__3255\
        );

    \I__402\ : InMux
    port map (
            O => \N__3267\,
            I => \N__3255\
        );

    \I__401\ : InMux
    port map (
            O => \N__3266\,
            I => \N__3255\
        );

    \I__400\ : InMux
    port map (
            O => \N__3265\,
            I => \N__3252\
        );

    \I__399\ : Odrv4
    port map (
            O => \N__3262\,
            I => \IR_ff7_q_ret_1_fast\
        );

    \I__398\ : LocalMux
    port map (
            O => \N__3255\,
            I => \IR_ff7_q_ret_1_fast\
        );

    \I__397\ : LocalMux
    port map (
            O => \N__3252\,
            I => \IR_ff7_q_ret_1_fast\
        );

    \I__396\ : CascadeMux
    port map (
            O => \N__3245\,
            I => \seq.counter.T_0_fast_RNIP4D21Z0Z_2_cascade_\
        );

    \I__395\ : CascadeMux
    port map (
            O => \N__3242\,
            I => \T_0_fast_RNILB791_2_cascade_\
        );

    \I__394\ : InMux
    port map (
            O => \N__3239\,
            I => \N__3236\
        );

    \I__393\ : LocalMux
    port map (
            O => \N__3236\,
            I => \N__3233\
        );

    \I__392\ : Span4Mux_s2_h
    port map (
            O => \N__3233\,
            I => \N__3230\
        );

    \I__391\ : Odrv4
    port map (
            O => \N__3230\,
            I => \pc.G_12_i_0\
        );

    \I__390\ : CascadeMux
    port map (
            O => \N__3227\,
            I => \seq.counter.T_0_fast_RNIG89VZ0Z_2_cascade_\
        );

    \I__389\ : InMux
    port map (
            O => \N__3224\,
            I => \N__3221\
        );

    \I__388\ : LocalMux
    port map (
            O => \N__3221\,
            I => \N__3218\
        );

    \I__387\ : Odrv4
    port map (
            O => \N__3218\,
            I => bus_6
        );

    \I__386\ : CascadeMux
    port map (
            O => \N__3215\,
            I => \N__3212\
        );

    \I__385\ : InMux
    port map (
            O => \N__3212\,
            I => \N__3207\
        );

    \I__384\ : InMux
    port map (
            O => \N__3211\,
            I => \N__3202\
        );

    \I__383\ : InMux
    port map (
            O => \N__3210\,
            I => \N__3202\
        );

    \I__382\ : LocalMux
    port map (
            O => \N__3207\,
            I => ir_out_fast_4
        );

    \I__381\ : LocalMux
    port map (
            O => \N__3202\,
            I => ir_out_fast_4
        );

    \I__380\ : CascadeMux
    port map (
            O => \N__3197\,
            I => \seq.counter.T_RNI0T6TZ0Z_4_cascade_\
        );

    \I__379\ : CascadeMux
    port map (
            O => \N__3194\,
            I => \N__3191\
        );

    \I__378\ : InMux
    port map (
            O => \N__3191\,
            I => \N__3188\
        );

    \I__377\ : LocalMux
    port map (
            O => \N__3188\,
            I => \N__3185\
        );

    \I__376\ : Span4Mux_s1_h
    port map (
            O => \N__3185\,
            I => \N__3177\
        );

    \I__375\ : InMux
    port map (
            O => \N__3184\,
            I => \N__3172\
        );

    \I__374\ : InMux
    port map (
            O => \N__3183\,
            I => \N__3172\
        );

    \I__373\ : InMux
    port map (
            O => \N__3182\,
            I => \N__3167\
        );

    \I__372\ : InMux
    port map (
            O => \N__3181\,
            I => \N__3167\
        );

    \I__371\ : InMux
    port map (
            O => \N__3180\,
            I => \N__3164\
        );

    \I__370\ : Odrv4
    port map (
            O => \N__3177\,
            I => ir_out_7_rep1
        );

    \I__369\ : LocalMux
    port map (
            O => \N__3172\,
            I => ir_out_7_rep1
        );

    \I__368\ : LocalMux
    port map (
            O => \N__3167\,
            I => ir_out_7_rep1
        );

    \I__367\ : LocalMux
    port map (
            O => \N__3164\,
            I => ir_out_7_rep1
        );

    \I__366\ : InMux
    port map (
            O => \N__3155\,
            I => \N__3148\
        );

    \I__365\ : InMux
    port map (
            O => \N__3154\,
            I => \N__3145\
        );

    \I__364\ : InMux
    port map (
            O => \N__3153\,
            I => \N__3140\
        );

    \I__363\ : InMux
    port map (
            O => \N__3152\,
            I => \N__3140\
        );

    \I__362\ : InMux
    port map (
            O => \N__3151\,
            I => \N__3137\
        );

    \I__361\ : LocalMux
    port map (
            O => \N__3148\,
            I => \N__3132\
        );

    \I__360\ : LocalMux
    port map (
            O => \N__3145\,
            I => \N__3132\
        );

    \I__359\ : LocalMux
    port map (
            O => \N__3140\,
            I => \N__3127\
        );

    \I__358\ : LocalMux
    port map (
            O => \N__3137\,
            I => \N__3127\
        );

    \I__357\ : Span4Mux_v
    port map (
            O => \N__3132\,
            I => \N__3124\
        );

    \I__356\ : Odrv12
    port map (
            O => \N__3127\,
            I => \seq_T_2_rep1\
        );

    \I__355\ : Odrv4
    port map (
            O => \N__3124\,
            I => \seq_T_2_rep1\
        );

    \I__354\ : CascadeMux
    port map (
            O => \N__3119\,
            I => \seq.D_1_0_x_cascade_\
        );

    \I__353\ : CascadeMux
    port map (
            O => \N__3116\,
            I => \ROM_OE_cascade_\
        );

    \I__352\ : InMux
    port map (
            O => \N__3113\,
            I => \N__3110\
        );

    \I__351\ : LocalMux
    port map (
            O => \N__3110\,
            I => \pc.program_counter_m_2\
        );

    \I__350\ : InMux
    port map (
            O => \N__3107\,
            I => \N__3103\
        );

    \I__349\ : InMux
    port map (
            O => \N__3106\,
            I => \N__3100\
        );

    \I__348\ : LocalMux
    port map (
            O => \N__3103\,
            I => \N__3097\
        );

    \I__347\ : LocalMux
    port map (
            O => \N__3100\,
            I => \pc.out_1_0_iv_0\
        );

    \I__346\ : Odrv12
    port map (
            O => \N__3097\,
            I => \pc.out_1_0_iv_0\
        );

    \I__345\ : CascadeMux
    port map (
            O => \N__3092\,
            I => \pc.G_10_0_a11_2_1_cascade_\
        );

    \I__344\ : InMux
    port map (
            O => \N__3089\,
            I => \N__3086\
        );

    \I__343\ : LocalMux
    port map (
            O => \N__3086\,
            I => \N__3083\
        );

    \I__342\ : Odrv4
    port map (
            O => \N__3083\,
            I => \pc.N_23\
        );

    \I__341\ : CascadeMux
    port map (
            O => \N__3080\,
            I => \pc.program_counter_RNO_6Z0Z_2_cascade_\
        );

    \I__340\ : InMux
    port map (
            O => \N__3077\,
            I => \N__3074\
        );

    \I__339\ : LocalMux
    port map (
            O => \N__3074\,
            I => \pc.G_10_0_a11_5_2\
        );

    \I__338\ : CascadeMux
    port map (
            O => \N__3071\,
            I => \seq.S1_1Z0Z_0_cascade_\
        );

    \I__337\ : CascadeMux
    port map (
            O => \N__3068\,
            I => \seq_S1_0_cascade_\
        );

    \I__336\ : InMux
    port map (
            O => \N__3065\,
            I => \N__3062\
        );

    \I__335\ : LocalMux
    port map (
            O => \N__3062\,
            I => \N__3059\
        );

    \I__334\ : Odrv4
    port map (
            O => \N__3059\,
            I => \pc.N_16\
        );

    \I__333\ : CascadeMux
    port map (
            O => \N__3056\,
            I => \ALU_main.N_48_cascade_\
        );

    \I__332\ : CascadeMux
    port map (
            O => \N__3053\,
            I => \alu_out_m_7_cascade_\
        );

    \I__331\ : CascadeMux
    port map (
            O => \N__3050\,
            I => \acc_out_m_7_cascade_\
        );

    \I__330\ : IoInMux
    port map (
            O => \N__3047\,
            I => \N__3044\
        );

    \I__329\ : LocalMux
    port map (
            O => \N__3044\,
            I => \N__3041\
        );

    \I__328\ : Span12Mux_s1_h
    port map (
            O => \N__3041\,
            I => \N__3038\
        );

    \I__327\ : Odrv12
    port map (
            O => \N__3038\,
            I => out_c_7
        );

    \I__326\ : InMux
    port map (
            O => \N__3035\,
            I => \N__3032\
        );

    \I__325\ : LocalMux
    port map (
            O => \N__3032\,
            I => \pc.out_1_2_iv_0\
        );

    \I__324\ : CascadeMux
    port map (
            O => \N__3029\,
            I => \pc.program_counter_RNO_7Z0Z_0_cascade_\
        );

    \I__323\ : InMux
    port map (
            O => \N__3026\,
            I => \N__3023\
        );

    \I__322\ : LocalMux
    port map (
            O => \N__3023\,
            I => \pc.program_counter_RNO_3Z0Z_0\
        );

    \I__321\ : InMux
    port map (
            O => \N__3020\,
            I => \N__3017\
        );

    \I__320\ : LocalMux
    port map (
            O => \N__3017\,
            I => \pc.program_counter_RNO_8Z0Z_0\
        );

    \I__319\ : CascadeMux
    port map (
            O => \N__3014\,
            I => \pc.program_counter_m_0_2_cascade_\
        );

    \I__318\ : CascadeMux
    port map (
            O => \N__3011\,
            I => \N__3008\
        );

    \I__317\ : InMux
    port map (
            O => \N__3008\,
            I => \N__3002\
        );

    \I__316\ : InMux
    port map (
            O => \N__3007\,
            I => \N__3002\
        );

    \I__315\ : LocalMux
    port map (
            O => \N__3002\,
            I => \AR_out_2\
        );

    \I__314\ : CascadeMux
    port map (
            O => \N__2999\,
            I => \N__2995\
        );

    \I__313\ : InMux
    port map (
            O => \N__2998\,
            I => \N__2992\
        );

    \I__312\ : InMux
    port map (
            O => \N__2995\,
            I => \N__2989\
        );

    \I__311\ : LocalMux
    port map (
            O => \N__2992\,
            I => \AR_out_0\
        );

    \I__310\ : LocalMux
    port map (
            O => \N__2989\,
            I => \AR_out_0\
        );

    \I__309\ : InMux
    port map (
            O => \N__2984\,
            I => \N__2981\
        );

    \I__308\ : LocalMux
    port map (
            O => \N__2981\,
            I => \mem_data_2_7_0__N_7_0\
        );

    \I__307\ : InMux
    port map (
            O => \N__2978\,
            I => \N__2975\
        );

    \I__306\ : LocalMux
    port map (
            O => \N__2975\,
            I => \pc.program_counter_m_0_0\
        );

    \I__305\ : CascadeMux
    port map (
            O => \N__2972\,
            I => \pc.out_1_2_iv_0_cascade_\
        );

    \I__304\ : CascadeMux
    port map (
            O => \N__2969\,
            I => \pc.tbuf.g0Z0Z_1_cascade_\
        );

    \I__303\ : InMux
    port map (
            O => \N__2966\,
            I => \N__2963\
        );

    \I__302\ : LocalMux
    port map (
            O => \N__2963\,
            I => bus_0
        );

    \I__301\ : InMux
    port map (
            O => \N__2960\,
            I => \N__2957\
        );

    \I__300\ : LocalMux
    port map (
            O => \N__2957\,
            I => \mem_data_2_7_0__N_14_0\
        );

    \I__299\ : CascadeMux
    port map (
            O => \N__2954\,
            I => \bus_6_cascade_\
        );

    \I__298\ : CascadeMux
    port map (
            O => \N__2951\,
            I => \N_5_0_cascade_\
        );

    \I__297\ : InMux
    port map (
            O => \N__2948\,
            I => \N__2945\
        );

    \I__296\ : LocalMux
    port map (
            O => \N__2945\,
            I => \N__2942\
        );

    \I__295\ : Span4Mux_v
    port map (
            O => \N__2942\,
            I => \N__2939\
        );

    \I__294\ : Odrv4
    port map (
            O => \N__2939\,
            I => \mem_data_2_7_0__g1\
        );

    \I__293\ : CascadeMux
    port map (
            O => \N__2936\,
            I => \seq_un1_IR_OE_4_1_cascade_\
        );

    \I__292\ : InMux
    port map (
            O => \N__2933\,
            I => \N__2930\
        );

    \I__291\ : LocalMux
    port map (
            O => \N__2930\,
            I => \N__2927\
        );

    \I__290\ : Span4Mux_h
    port map (
            O => \N__2927\,
            I => \N__2924\
        );

    \I__289\ : Odrv4
    port map (
            O => \N__2924\,
            I => \pc.program_counter_RNO_5Z0Z_0\
        );

    \I__288\ : CascadeMux
    port map (
            O => \N__2921\,
            I => \seq.un17_IR_OE_cascade_\
        );

    \I__287\ : CascadeMux
    port map (
            O => \N__2918\,
            I => \seq_PC_LD_0_0_cascade_\
        );

    \I__286\ : InMux
    port map (
            O => \N__2915\,
            I => \N__2912\
        );

    \I__285\ : LocalMux
    port map (
            O => \N__2912\,
            I => \seq.D_6_x\
        );

    \I__284\ : CascadeMux
    port map (
            O => \N__2909\,
            I => \pc.program_counter_m_3_cascade_\
        );

    \I__283\ : InMux
    port map (
            O => \N__2906\,
            I => \N__2903\
        );

    \I__282\ : LocalMux
    port map (
            O => \N__2903\,
            I => \pc.tbuf.gZ0Z3\
        );

    \I__281\ : CascadeMux
    port map (
            O => \N__2900\,
            I => \pc.tbuf.g0Z0Z_3_cascade_\
        );

    \I__280\ : CascadeMux
    port map (
            O => \N__2897\,
            I => \bus_3_cascade_\
        );

    \I__279\ : CascadeMux
    port map (
            O => \N__2894\,
            I => \N__2891\
        );

    \I__278\ : InMux
    port map (
            O => \N__2891\,
            I => \N__2888\
        );

    \I__277\ : LocalMux
    port map (
            O => \N__2888\,
            I => \N__2885\
        );

    \I__276\ : Odrv4
    port map (
            O => \N__2885\,
            I => \seq_MAR_LD_1_0\
        );

    \I__275\ : CascadeMux
    port map (
            O => \N__2882\,
            I => \N__2879\
        );

    \I__274\ : InMux
    port map (
            O => \N__2879\,
            I => \N__2876\
        );

    \I__273\ : LocalMux
    port map (
            O => \N__2876\,
            I => \pc.program_counter_m_3\
        );

    \I__272\ : CascadeMux
    port map (
            O => \N__2873\,
            I => \seq.DZ0Z_0_cascade_\
        );

    \I__271\ : InMux
    port map (
            O => \N__2870\,
            I => \N__2867\
        );

    \I__270\ : LocalMux
    port map (
            O => \N__2867\,
            I => clk_c
        );

    \I__269\ : IoInMux
    port map (
            O => \N__2864\,
            I => \N__2861\
        );

    \I__268\ : LocalMux
    port map (
            O => \N__2861\,
            I => buf_clk_1
        );

    \I__267\ : CascadeMux
    port map (
            O => \N__2858\,
            I => \pc.N_21_0_cascade_\
        );

    \I__266\ : CascadeMux
    port map (
            O => \N__2855\,
            I => \seq_D_6_cascade_\
        );

    \I__265\ : InMux
    port map (
            O => \N__2852\,
            I => \N__2849\
        );

    \I__264\ : LocalMux
    port map (
            O => \N__2849\,
            I => \pc.G_12_i_a3_1\
        );

    \INVout_reg.ff4.qC\ : INV
    port map (
            O => \INVout_reg.ff4.qC_net\,
            I => \N__4804\
        );

    \INVb_reg.ff4.qC\ : INV
    port map (
            O => \INVb_reg.ff4.qC_net\,
            I => \N__4807\
        );

    \INVout_reg.ff2.qC\ : INV
    port map (
            O => \INVout_reg.ff2.qC_net\,
            I => \N__4803\
        );

    \INVb_reg.ff3.qC\ : INV
    port map (
            O => \INVb_reg.ff3.qC_net\,
            I => \N__4799\
        );

    \INVIR.ff1.q_nerC\ : INV
    port map (
            O => \INVIR.ff1.q_nerC_net\,
            I => \N__4795\
        );

    \INVout_reg.ff3.qC\ : INV
    port map (
            O => \INVout_reg.ff3.qC_net\,
            I => \N__4788\
        );

    \INVout_reg.ff6.qC\ : INV
    port map (
            O => \INVout_reg.ff6.qC_net\,
            I => \N__4808\
        );

    \INVb_reg.ff2.qC\ : INV
    port map (
            O => \INVb_reg.ff2.qC_net\,
            I => \N__4806\
        );

    \INVout_reg.ff7.qC\ : INV
    port map (
            O => \INVout_reg.ff7.qC_net\,
            I => \N__4802\
        );

    \INVb_reg.ff6.qC\ : INV
    port map (
            O => \INVb_reg.ff6.qC_net\,
            I => \N__4798\
        );

    \INVmar.ff4.q_nerC\ : INV
    port map (
            O => \INVmar.ff4.q_nerC_net\,
            I => \N__4794\
        );

    \INVacc.ff1.qC\ : INV
    port map (
            O => \INVacc.ff1.qC_net\,
            I => \N__4791\
        );

    \INVIR.ff2.q_nerC\ : INV
    port map (
            O => \INVIR.ff2.q_nerC_net\,
            I => \N__4783\
        );

    \INVacc.ff7.qC\ : INV
    port map (
            O => \INVacc.ff7.qC_net\,
            I => \N__4801\
        );

    \INVb_reg.ff5.qC\ : INV
    port map (
            O => \INVb_reg.ff5.qC_net\,
            I => \N__4797\
        );

    \INVAR.ff2.qC\ : INV
    port map (
            O => \INVAR.ff2.qC_net\,
            I => \N__4779\
        );

    \INVseq.q_retC\ : INV
    port map (
            O => \INVseq.q_retC_net\,
            I => \N__4805\
        );

    \INVseq.q_ret_1C\ : INV
    port map (
            O => \INVseq.q_ret_1C_net\,
            I => \N__4800\
        );

    \INVseq.counter.T_0C\ : INV
    port map (
            O => \INVseq.counter.T_0C_net\,
            I => \N__4782\
        );

    \INVIR.ff7.q_0_nerC\ : INV
    port map (
            O => \INVIR.ff7.q_0_nerC_net\,
            I => \N__4793\
        );

    \INVseq.counter.T_0_fast_2C\ : INV
    port map (
            O => \INVseq.counter.T_0_fast_2C_net\,
            I => \N__4790\
        );

    \INVIR.ff6.q_ret_1C\ : INV
    port map (
            O => \INVIR.ff6.q_ret_1C_net\,
            I => \N__4785\
        );

    \INVIR.ff7.q_0_fastC\ : INV
    port map (
            O => \INVIR.ff7.q_0_fastC_net\,
            I => \N__4781\
        );

    \INVmar.ff1.q_nerC\ : INV
    port map (
            O => \INVmar.ff1.q_nerC_net\,
            I => \N__4778\
        );

    \INVout_reg.ff8.qC\ : INV
    port map (
            O => \INVout_reg.ff8.qC_net\,
            I => \N__4776\
        );

    \INVAR.ff3.qC\ : INV
    port map (
            O => \INVAR.ff3.qC_net\,
            I => \N__4777\
        );

    \INVseq.counter.T_4C\ : INV
    port map (
            O => \INVseq.counter.T_4C_net\,
            I => \N__4792\
        );

    \INVIR.ff5.q_0_nerC\ : INV
    port map (
            O => \INVIR.ff5.q_0_nerC_net\,
            I => \N__4789\
        );

    \INVIR.ff7.q_ret_1C\ : INV
    port map (
            O => \INVIR.ff7.q_ret_1C_net\,
            I => \N__4784\
        );

    \INVIR.ff5.q_0_rep1C\ : INV
    port map (
            O => \INVIR.ff5.q_0_rep1C_net\,
            I => \N__4780\
        );

    \INVAR.ff4.qC\ : INV
    port map (
            O => \INVAR.ff4.qC_net\,
            I => \N__4775\
        );

    \INVseq.counter.T_0_2_rep1C\ : INV
    port map (
            O => \INVseq.counter.T_0_2_rep1C_net\,
            I => \N__4774\
        );

    \IN_MUX_bfv_4_12_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "00"
        )
    port map (
            carryinitin => '0',
            carryinitout => \bfn_4_12_0_\
        );

    \IN_MUX_bfv_4_13_0_\ : ICE_CARRY_IN_MUX
    generic map (
            C_INIT => "10"
        )
    port map (
            carryinitin => \ALU_main.un1_A_cry_6\,
            carryinitout => \bfn_4_13_0_\
        );

    \buf_clk_1_inferred_clock_0_RNIEA29\ : ICE_GB
    port map (
            USERSIGNALTOGLOBALBUFFER => \N__2864\,
            GLOBALBUFFEROUTPUT => buf_clk_1_g
        );

    \GND\ : GND
    port map (
            Y => \GNDG0\
        );

    \VCC\ : VCC
    port map (
            Y => \VCCG0\
        );

    \GND_Inst\ : GND
    port map (
            Y => \_gnd_net_\
        );

    \seq.counter.T_0_2_rep1_LC_1_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010101010101010"
        )
    port map (
            in0 => \N__8666\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \_gnd_net_\,
            lcout => \seq_T_2_rep1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVseq.counter.T_0_2_rep1C_net\,
            ce => 'H',
            sr => \N__7288\
        );

    \AR.ff1.q_LC_1_8_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110110001001100"
        )
    port map (
            in0 => \N__4273\,
            in1 => \N__2998\,
            in2 => \N__4668\,
            in3 => \N__2966\,
            lcout => \AR_out_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVseq.counter.T_0_2_rep1C_net\,
            ce => 'H',
            sr => \N__7288\
        );

    \seq.counter.T_0_2_LC_1_8_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8665\,
            lcout => \seq_T_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVseq.counter.T_0_2_rep1C_net\,
            ce => 'H',
            sr => \N__7288\
        );

    \buf_clk_1_inferred_clock_0_RNO_LC_1_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100000000"
        )
    port map (
            in0 => \N__4337\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__2870\,
            lcout => buf_clk_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNI1BHH1_0_LC_1_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__3643\,
            in1 => \N__4639\,
            in2 => \N__3548\,
            in3 => \N__4252\,
            lcout => \pc.program_counter_m_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_4_0_LC_1_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001010100000000"
        )
    port map (
            in0 => \N__3541\,
            in1 => \N__4251\,
            in2 => \N__4654\,
            in3 => \N__4205\,
            lcout => OPEN,
            ltout => \pc.N_21_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_1_0_LC_1_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101000100000000"
        )
    port map (
            in0 => \N__8672\,
            in1 => \N__3644\,
            in2 => \N__2858\,
            in3 => \N__2933\,
            lcout => \pc.G_12_i_a3_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mar.ff1.q_sbtinv_LC_1_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010111011111111"
        )
    port map (
            in0 => \N__3545\,
            in1 => \N__4640\,
            in2 => \N__2894\,
            in3 => \N__4497\,
            lcout => \mar.MAR_LD_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_10_2_LC_1_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__3718\,
            in1 => \N__3152\,
            in2 => \N__3537\,
            in3 => \N__4248\,
            lcout => \pc.program_counter_m_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.decoder.D_6_LC_1_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__5455\,
            in1 => \N__3302\,
            in2 => \N__3194\,
            in3 => \N__5408\,
            lcout => \seq_D_6\,
            ltout => \seq_D_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNI0GCL1_1_LC_1_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__3523\,
            in1 => \N__4837\,
            in2 => \N__2855\,
            in3 => \N__3153\,
            lcout => \pc.program_counter_m_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_0_LC_1_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000101010101"
        )
    port map (
            in0 => \N__3239\,
            in1 => \N__2852\,
            in2 => \N__3590\,
            in3 => \N__3026\,
            lcout => \pc.program_counterZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4773\,
            ce => 'H',
            sr => \N__7287\
        );

    \pc.tbuf.g3_LC_1_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001110111"
        )
    port map (
            in0 => \N__2948\,
            in1 => \N__7121\,
            in2 => \_gnd_net_\,
            in3 => \N__6482\,
            lcout => \pc.tbuf.gZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNI2ICL1_3_LC_1_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010100010100000"
        )
    port map (
            in0 => \N__4009\,
            in1 => \N__4249\,
            in2 => \N__3547\,
            in3 => \N__3155\,
            lcout => \pc.program_counter_m_3\,
            ltout => \pc.program_counter_m_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.tbuf.g0_3_LC_1_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__4485\,
            in1 => \N__3890\,
            in2 => \N__2909\,
            in3 => \N__2906\,
            lcout => \pc.tbuf.g0Z0Z_3\,
            ltout => \pc.tbuf.g0Z0Z_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.tbuf.g0_LC_1_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111111101"
        )
    port map (
            in0 => \N__7618\,
            in1 => \N__7749\,
            in2 => \N__2900\,
            in3 => \N__7544\,
            lcout => OPEN,
            ltout => \bus_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \AR.ff4.q_LC_1_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110010011001100"
        )
    port map (
            in0 => \N__4250\,
            in1 => \N__3912\,
            in2 => \N__2897\,
            in3 => \N__4669\,
            lcout => \AR.ff4.AR_out_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVAR.ff4.qC_net\,
            ce => 'H',
            sr => \N__7289\
        );

    \seq.MAR_LD_1_0_LC_1_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4965\,
            in1 => \N__5138\,
            in2 => \_gnd_net_\,
            in3 => \N__5005\,
            lcout => \seq_MAR_LD_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.g2_0_LC_1_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000101"
        )
    port map (
            in0 => \N__5004\,
            in1 => \_gnd_net_\,
            in2 => \N__5147\,
            in3 => \N__4964\,
            lcout => \seq.g2Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.tbuf.out_1_iv_1_1_LC_1_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101100000011"
        )
    port map (
            in0 => \N__3328\,
            in1 => \N__3888\,
            in2 => \N__2882\,
            in3 => \N__4541\,
            lcout => \pc.out_1_iv_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.decoder.D_0_LC_1_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__3434\,
            in1 => \N__3272\,
            in2 => \N__3215\,
            in3 => \N__5500\,
            lcout => \seq.DZ0Z_0\,
            ltout => \seq.DZ0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_0_2_rep1_RNIE27K3_LC_1_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101010111"
        )
    port map (
            in0 => \N__3151\,
            in1 => \N__5134\,
            in2 => \N__2873\,
            in3 => \N__5003\,
            lcout => \seq_un1_IR_OE_4_1\,
            ltout => \seq_un1_IR_OE_4_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_3_2_LC_1_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111101010101"
        )
    port map (
            in0 => \N__4539\,
            in1 => \N__4457\,
            in2 => \N__2936\,
            in3 => \N__4194\,
            lcout => \pc.G_10_0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_5_0_LC_1_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111100001111"
        )
    port map (
            in0 => \N__4540\,
            in1 => \N__3327\,
            in2 => \N__8765\,
            in3 => \N__4458\,
            lcout => \pc.program_counter_RNO_5Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_8_2_LC_1_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__8667\,
            in1 => \N__4547\,
            in2 => \N__3722\,
            in3 => \N__4183\,
            lcout => \pc.N_23\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.q_ret_RNI7NFN_LC_1_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100000000000000"
        )
    port map (
            in0 => \N__3184\,
            in1 => \N__5561\,
            in2 => \N__4292\,
            in3 => \N__5398\,
            lcout => OPEN,
            ltout => \seq.un17_IR_OE_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_RNIPKHM1_3_LC_1_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100001111"
        )
    port map (
            in0 => \N__5218\,
            in1 => \N__2915\,
            in2 => \N__2921\,
            in3 => \N__3301\,
            lcout => \seq_PC_LD_0_0\,
            ltout => \seq_PC_LD_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_0_3_LC_1_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110011101111"
        )
    port map (
            in0 => \N__4184\,
            in1 => \N__3560\,
            in2 => \N__2918\,
            in3 => \N__8668\,
            lcout => \pc.g0_rn_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.decoder.D_6_x_LC_1_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000100010"
        )
    port map (
            in0 => \N__5397\,
            in1 => \N__5443\,
            in2 => \_gnd_net_\,
            in3 => \N__3183\,
            lcout => \seq.D_6_x\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \IR.ff5.q_0_rep1_LC_1_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101000001010"
        )
    port map (
            in0 => \N__5562\,
            in1 => \_gnd_net_\,
            in2 => \N__8686\,
            in3 => \N__5594\,
            lcout => ir_out_4_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVIR.ff5.q_0_rep1C_net\,
            ce => 'H',
            sr => \N__7294\
        );

    \seq.decoder.D_4_0_LC_1_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001000000"
        )
    port map (
            in0 => \N__5444\,
            in1 => \N__5494\,
            in2 => \N__5407\,
            in3 => \N__3180\,
            lcout => \seq.D_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf1.out_1_0_iv_LC_1_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__6829\,
            in1 => \N__6789\,
            in2 => \N__6746\,
            in3 => \N__6521\,
            lcout => bus_6,
            ltout => \bus_6_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \IR.ff7.q_0_ner_RNI7C4KI_LC_1_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8660\,
            in2 => \N__2954\,
            in3 => \N__3964\,
            lcout => \N_5_0\,
            ltout => \N_5_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \IR.ff7.q_ret_1_LC_1_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000111100001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__2951\,
            in3 => \_gnd_net_\,
            lcout => ir_out_i_2_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVIR.ff7.q_ret_1C_net\,
            ce => 'H',
            sr => \N__7298\
        );

    \seq.g0_i_a3_2_LC_1_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010000000000"
        )
    port map (
            in0 => \N__5545\,
            in1 => \N__3295\,
            in2 => \_gnd_net_\,
            in3 => \N__3374\,
            lcout => \seq.g0_i_a3Z0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \IR.ff6.q_0_fast_LC_1_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8661\,
            in1 => \N__6086\,
            in2 => \_gnd_net_\,
            in3 => \N__4417\,
            lcout => \IR_ff6_q_0_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVIR.ff7.q_ret_1C_net\,
            ce => 'H',
            sr => \N__7298\
        );

    \seq.decoder.D_3_0_LC_1_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__5445\,
            in1 => \N__3296\,
            in2 => \N__3424\,
            in3 => \N__3265\,
            lcout => \seq.D_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \IR.ff7.q_ret_1_fast_LC_1_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4351\,
            lcout => \IR_ff7_q_ret_1_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVIR.ff7.q_ret_1C_net\,
            ce => 'H',
            sr => \N__7298\
        );

    \IR.ff5.q_0_ner_LC_1_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__7995\,
            in1 => \N__7964\,
            in2 => \N__7922\,
            in3 => \N__7388\,
            lcout => ir_out_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVIR.ff5.q_0_nerC_net\,
            ce => \N__8683\,
            sr => \N__7303\
        );

    \seq.counter.T_4_LC_1_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5222\,
            lcout => \seq.counter.TZ0Z_4\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVseq.counter.T_4C_net\,
            ce => 'H',
            sr => \N__7306\
        );

    \mem.data_2_7_0__g1_LC_2_7_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011101110"
        )
    port map (
            in0 => \N__7044\,
            in1 => \N__7186\,
            in2 => \_gnd_net_\,
            in3 => \N__6965\,
            lcout => \mem_data_2_7_0__g1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.tbuf.out_1_0_iv_0_LC_2_8_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111100010001000"
        )
    port map (
            in0 => \N__3007\,
            in1 => \N__4204\,
            in2 => \N__5993\,
            in3 => \N__7441\,
            lcout => \pc.out_1_0_iv_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNI3DHH1_2_LC_2_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100100010001000"
        )
    port map (
            in0 => \N__3546\,
            in1 => \N__3711\,
            in2 => \N__4666\,
            in3 => \N__4271\,
            lcout => OPEN,
            ltout => \pc.program_counter_m_0_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.tbuf.g0_9_LC_2_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111101"
        )
    port map (
            in0 => \N__2960\,
            in1 => \N__3106\,
            in2 => \N__3014\,
            in3 => \N__6522\,
            lcout => \pc.tbuf.g0_1_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \AR.ff3.q_LC_2_8_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111100001110000"
        )
    port map (
            in0 => \N__4272\,
            in1 => \N__4644\,
            in2 => \N__3011\,
            in3 => \N__3455\,
            lcout => \AR_out_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVAR.ff3.qC_net\,
            ce => 'H',
            sr => \N__7291\
        );

    \mem.data_2_7_0__g0_2_LC_2_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110110101"
        )
    port map (
            in0 => \N__7130\,
            in1 => \N__7057\,
            in2 => \N__7196\,
            in3 => \N__6967\,
            lcout => \mem_data_2_7_0__N_7_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.tbuf.out_1_2_iv_0_LC_2_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__6067\,
            in1 => \N__4203\,
            in2 => \N__2999\,
            in3 => \N__7398\,
            lcout => \pc.out_1_2_iv_0\,
            ltout => \pc.out_1_2_iv_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.tbuf.g0_5_LC_2_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111110011111101"
        )
    port map (
            in0 => \N__2984\,
            in1 => \N__2978\,
            in2 => \N__2972\,
            in3 => \N__6523\,
            lcout => \pc.tbuf.g0Z0Z_1\,
            ltout => \pc.tbuf.g0Z0Z_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.tbuf.g0_4_LC_2_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110100"
        )
    port map (
            in0 => \N__8877\,
            in1 => \N__8764\,
            in2 => \N__2969\,
            in3 => \N__8814\,
            lcout => bus_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mem.data_2_7_0__g0_3_LC_2_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110100111"
        )
    port map (
            in0 => \N__6966\,
            in1 => \N__7192\,
            in2 => \N__7058\,
            in3 => \N__7129\,
            lcout => \mem_data_2_7_0__N_14_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.ALU_Out_0_7_LC_2_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001100110"
        )
    port map (
            in0 => \N__6269\,
            in1 => \N__5875\,
            in2 => \_gnd_net_\,
            in3 => \N__6194\,
            lcout => OPEN,
            ltout => \ALU_main.N_48_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.un1_A_cry_6_c_RNIGN9C9_LC_2_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__3791\,
            in1 => \N__5742\,
            in2 => \N__3056\,
            in3 => \N__5644\,
            lcout => alu_out_m_7,
            ltout => \alu_out_m_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf1.out_1_iv_LC_2_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111110001"
        )
    port map (
            in0 => \N__6465\,
            in1 => \N__6901\,
            in2 => \N__3053\,
            in3 => \N__6327\,
            lcout => bus_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acc.ff8.q_RNI449H1_LC_2_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5876\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7399\,
            lcout => acc_out_m_7,
            ltout => \acc_out_m_7_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \out_reg.ff8.q_LC_2_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111110011111101"
        )
    port map (
            in0 => \N__6466\,
            in1 => \N__6293\,
            in2 => \N__3050\,
            in3 => \N__6902\,
            lcout => out_c_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVout_reg.ff8.qC_net\,
            ce => \N__7480\,
            sr => \N__7290\
        );

    \pc.program_counter_RNO_7_0_LC_2_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100100010"
        )
    port map (
            in0 => \N__6221\,
            in1 => \N__3035\,
            in2 => \_gnd_net_\,
            in3 => \N__6464\,
            lcout => OPEN,
            ltout => \pc.program_counter_RNO_7Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_3_0_LC_2_10_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000001010000"
        )
    port map (
            in0 => \N__3065\,
            in1 => \N__3020\,
            in2 => \N__3029\,
            in3 => \N__5033\,
            lcout => \pc.program_counter_RNO_3Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_8_0_LC_2_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5741\,
            in2 => \_gnd_net_\,
            in3 => \N__5643\,
            lcout => \pc.program_counter_RNO_8Z0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mem.data_2_7_0__g0_LC_2_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100100011001000"
        )
    port map (
            in0 => \N__7174\,
            in1 => \N__7118\,
            in2 => \N__7043\,
            in3 => \N__6933\,
            lcout => \mem_data_2_7_0__N_16_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mar.ff1.q_ner_LC_2_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__8908\,
            in1 => \N__8763\,
            in2 => \N__8878\,
            in3 => \N__8807\,
            lcout => mar_out_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVmar.ff1.q_nerC_net\,
            ce => \N__6382\,
            sr => \N__7292\
        );

    \seq.counter.T_RNI4RN46_3_LC_2_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000011100000000"
        )
    port map (
            in0 => \N__5217\,
            in1 => \N__4963\,
            in2 => \N__8684\,
            in3 => \N__3311\,
            lcout => \ROM_OE\,
            ltout => \ROM_OE_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_7_2_LC_2_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000100"
        )
    port map (
            in0 => \N__6934\,
            in1 => \N__7018\,
            in2 => \N__3116\,
            in3 => \N__7120\,
            lcout => \pc.G_10_0_a11_5_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_9_2_LC_2_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000001000000000"
        )
    port map (
            in0 => \N__7173\,
            in1 => \N__7119\,
            in2 => \N__7042\,
            in3 => \N__6932\,
            lcout => OPEN,
            ltout => \pc.G_10_0_a11_2_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_6_2_LC_2_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011111110"
        )
    port map (
            in0 => \N__3113\,
            in1 => \N__3107\,
            in2 => \N__3092\,
            in3 => \N__6463\,
            lcout => OPEN,
            ltout => \pc.program_counter_RNO_6Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_2_2_LC_2_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101010"
        )
    port map (
            in0 => \N__3089\,
            in1 => \N__3769\,
            in2 => \N__3080\,
            in3 => \N__3077\,
            lcout => \pc.G_10_0_sx\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.S1_1_0_LC_2_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__5499\,
            in1 => \N__3211\,
            in2 => \_gnd_net_\,
            in3 => \N__5405\,
            lcout => OPEN,
            ltout => \seq.S1_1Z0Z_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_RNIMQC72_4_LC_2_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010111011111"
        )
    port map (
            in0 => \N__5350\,
            in1 => \N__3182\,
            in2 => \N__3071\,
            in3 => \N__4897\,
            lcout => \seq_S1_0\,
            ltout => \seq_S1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_9_0_LC_2_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100100000010"
        )
    port map (
            in0 => \N__6245\,
            in1 => \N__6186\,
            in2 => \N__3068\,
            in3 => \N__6068\,
            lcout => \pc.N_16\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \IR.ff7.q_0_fast_LC_2_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1100110010101010"
        )
    port map (
            in0 => \N__3967\,
            in1 => \N__3224\,
            in2 => \_gnd_net_\,
            in3 => \N__8663\,
            lcout => \IR_ff7_q_0_fast\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVIR.ff7.q_0_fastC_net\,
            ce => 'H',
            sr => \N__7295\
        );

    \IR.ff5.q_0_fast_LC_2_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__5590\,
            in1 => \N__8662\,
            in2 => \_gnd_net_\,
            in3 => \N__5564\,
            lcout => ir_out_fast_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVIR.ff7.q_0_fastC_net\,
            ce => 'H',
            sr => \N__7295\
        );

    \seq.counter.T_RNI0T6T_4_LC_2_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__3210\,
            in1 => \N__3181\,
            in2 => \N__5362\,
            in3 => \N__5498\,
            lcout => OPEN,
            ltout => \seq.counter.T_RNI0T6TZ0Z_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_RNI0TT62_4_LC_2_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__3476\,
            in1 => \N__3966\,
            in2 => \N__3197\,
            in3 => \N__3386\,
            lcout => \seq_S0_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \IR.ff8.q_0_rep1_LC_2_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1011101110001000"
        )
    port map (
            in0 => \N__4383\,
            in1 => \N__8664\,
            in2 => \_gnd_net_\,
            in3 => \N__5311\,
            lcout => ir_out_7_rep1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVIR.ff7.q_0_fastC_net\,
            ce => 'H',
            sr => \N__7295\
        );

    \seq.decoder.D_1_0_x_LC_2_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__5497\,
            in1 => \N__3428\,
            in2 => \_gnd_net_\,
            in3 => \N__3268\,
            lcout => OPEN,
            ltout => \seq.D_1_0_x_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_0_2_rep1_RNIC9OP2_LC_2_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011011101110111"
        )
    port map (
            in0 => \N__4890\,
            in1 => \N__3154\,
            in2 => \N__3119\,
            in3 => \N__5448\,
            lcout => \seq_MAR_LD_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \IR.ff6.q_ret_1_LC_2_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0000000011111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4316\,
            lcout => ir_out_i_2_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVIR.ff6.q_ret_1C_net\,
            ce => 'H',
            sr => \N__7299\
        );

    \seq.B_LD_2_tz_LC_2_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000110011"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4889\,
            in2 => \_gnd_net_\,
            in3 => \N__5002\,
            lcout => \seq.B_LD_0_2_tz\,
            ltout => \seq.B_LD_0_2_tz_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_RNIR83I4_0_3_LC_2_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010101110101"
        )
    port map (
            in0 => \N__5216\,
            in1 => \N__5133\,
            in2 => \N__3314\,
            in3 => \N__5078\,
            lcout => \seq.counter.T_RNIR83I4_0Z0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.decoder.D_2_0_LC_2_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010000000000"
        )
    port map (
            in0 => \N__5446\,
            in1 => \N__3267\,
            in2 => \N__3432\,
            in3 => \N__3297\,
            lcout => \seq.D_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.decoder.D_1_0_LC_2_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000100000000000"
        )
    port map (
            in0 => \N__3266\,
            in1 => \N__5496\,
            in2 => \N__3433\,
            in3 => \N__5447\,
            lcout => \seq.D_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_RNIGQT43_1_LC_2_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100010001"
        )
    port map (
            in0 => \N__4542\,
            in1 => \N__8654\,
            in2 => \_gnd_net_\,
            in3 => \N__4179\,
            lcout => \N_30\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_0_fast_RNIP4D21_2_LC_2_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__3351\,
            in1 => \N__4413\,
            in2 => \N__3965\,
            in3 => \N__5290\,
            lcout => OPEN,
            ltout => \seq.counter.T_0_fast_RNIP4D21Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_0_fast_RNILB791_2_LC_2_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000010101010"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3245\,
            in3 => \N__5548\,
            lcout => \T_0_fast_RNILB791_2\,
            ltout => \T_0_fast_RNILB791_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_0_0_LC_2_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100110001000"
        )
    port map (
            in0 => \N__8655\,
            in1 => \N__3671\,
            in2 => \N__3242\,
            in3 => \N__4543\,
            lcout => \pc.G_12_i_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_0_fast_2_LC_2_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__8659\,
            lcout => \seq.counter.T_fast_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVseq.counter.T_0_fast_2C_net\,
            ce => 'H',
            sr => \N__7304\
        );

    \seq.counter.T_0_fast_RNIG89V_2_LC_2_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000000000000000"
        )
    port map (
            in0 => \N__3377\,
            in1 => \N__3409\,
            in2 => \N__3355\,
            in3 => \N__5495\,
            lcout => OPEN,
            ltout => \seq.counter.T_0_fast_RNIG89VZ0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_0_fast_RNICF361_2_LC_2_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101011110000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__3227\,
            in3 => \N__5549\,
            lcout => \OUT_LD\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \IR.ff8.q_0_fast_LC_2_14_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1010111110100000"
        )
    port map (
            in0 => \N__4387\,
            in1 => \_gnd_net_\,
            in2 => \N__8685\,
            in3 => \N__5291\,
            lcout => ir_out_fast_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVseq.counter.T_0_fast_2C_net\,
            ce => 'H',
            sr => \N__7304\
        );

    \IR.ff7.q_0_ner_LC_2_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110001"
        )
    port map (
            in0 => \N__6525\,
            in1 => \N__6745\,
            in2 => \N__6836\,
            in3 => \N__6791\,
            lcout => ir_out_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVIR.ff7.q_0_nerC_net\,
            ce => \N__8687\,
            sr => \N__7307\
        );

    \IR.ff6.q_0_ner_LC_2_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__6692\,
            in1 => \N__6641\,
            in2 => \N__6605\,
            in3 => \N__6524\,
            lcout => ir_out_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVIR.ff7.q_0_nerC_net\,
            ce => \N__8687\,
            sr => \N__7307\
        );

    \IR.ff8.q_0_ner_LC_2_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111110001"
        )
    port map (
            in0 => \N__6526\,
            in1 => \N__6900\,
            in2 => \N__6309\,
            in3 => \N__6334\,
            lcout => ir_out_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVIR.ff7.q_0_nerC_net\,
            ce => \N__8687\,
            sr => \N__7307\
        );

    \seq.S0_0_i_N_3L3_LC_2_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5281\,
            in2 => \_gnd_net_\,
            in3 => \N__3375\,
            lcout => \seq.S0_0_i_N_3LZ0Z3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.un1_ALU_en_0_1_LC_2_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000101000001010"
        )
    port map (
            in0 => \N__3376\,
            in1 => \_gnd_net_\,
            in2 => \N__5299\,
            in3 => \_gnd_net_\,
            lcout => \seq.un1_ALU_en_0Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \IR.ff4.q_ner_LC_2_15_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__7740\,
            in1 => \N__7681\,
            in2 => \N__7593\,
            in3 => \N__7545\,
            lcout => ir_out_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVIR.ff7.q_0_nerC_net\,
            ce => \N__8687\,
            sr => \N__7307\
        );

    \seq.counter.T_0_fast_RNIOL5V_2_LC_2_16_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100000000000"
        )
    port map (
            in0 => \N__3356\,
            in1 => \N__4412\,
            in2 => \_gnd_net_\,
            in3 => \N__5547\,
            lcout => \seq_un1_AR_OE_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.tbuf.g2_LC_2_16_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110101010101"
        )
    port map (
            in0 => \N__3875\,
            in1 => \N__3335\,
            in2 => \_gnd_net_\,
            in3 => \N__4587\,
            lcout => \pc.tbuf.gZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \AR.ff4.q_RNIT1RE_LC_2_16_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__3963\,
            in1 => \N__3926\,
            in2 => \_gnd_net_\,
            in3 => \N__5295\,
            lcout => OPEN,
            ltout => \g0_0_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.tbuf.g0_1_LC_2_16_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110110010100000"
        )
    port map (
            in0 => \N__3985\,
            in1 => \N__5827\,
            in2 => \N__3479\,
            in3 => \N__7400\,
            lcout => \pc.tbuf.g0_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_RNIUILR_4_LC_2_16_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010001000"
        )
    port map (
            in0 => \N__5325\,
            in1 => \N__4411\,
            in2 => \_gnd_net_\,
            in3 => \N__5546\,
            lcout => \seq.counter.un7_ACC_LD_0\,
            ltout => \seq.counter.un7_ACC_LD_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_RNIK9TB2_4_LC_2_16_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__3467\,
            in1 => \N__5326\,
            in2 => \N__3461\,
            in3 => \N__5088\,
            lcout => \seq_un1_ALU_en_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_0_RNILSL08_1_2_LC_4_8_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000000000"
        )
    port map (
            in0 => \N__4667\,
            in1 => \N__4589\,
            in2 => \N__4943\,
            in3 => \N__4502\,
            lcout => \IR_OE_2\,
            ltout => \IR_OE_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.tbuf.g0_8_LC_4_8_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__8435\,
            in1 => \N__8448\,
            in2 => \N__3458\,
            in3 => \N__8279\,
            lcout => bus_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_0_1_LC_4_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111101111000"
        )
    port map (
            in0 => \N__3670\,
            in1 => \N__8553\,
            in2 => \N__4838\,
            in3 => \N__3599\,
            lcout => \pc.program_counter_4_rn_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.un1_inc_LC_4_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__8552\,
            in1 => \N__4578\,
            in2 => \_gnd_net_\,
            in3 => \N__4213\,
            lcout => \pc.un1_inc_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_4_3_LC_4_9_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3704\,
            in2 => \_gnd_net_\,
            in3 => \N__4832\,
            lcout => \pc.g1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_0_RNILSL08_2_LC_4_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000110000000000"
        )
    port map (
            in0 => \N__3446\,
            in1 => \N__4577\,
            in2 => \N__4686\,
            in3 => \N__4492\,
            lcout => \IR_OE_1\,
            ltout => \IR_OE_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_1_1_LC_4_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8114\,
            in2 => \N__3602\,
            in3 => \N__3598\,
            lcout => \pc.program_counter_4_sn_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_RNIAFFM9_4_LC_4_9_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101110000001100"
        )
    port map (
            in0 => \N__5761\,
            in1 => \N__3731\,
            in2 => \N__5684\,
            in3 => \N__3824\,
            lcout => alu_out_m_0_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_2_0_LC_4_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000010001000100"
        )
    port map (
            in0 => \N__4580\,
            in1 => \N__3578\,
            in2 => \N__4694\,
            in3 => \N__4267\,
            lcout => \pc.G_12_i_a3_2_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_6_0_LC_4_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__8549\,
            in1 => \N__8756\,
            in2 => \_gnd_net_\,
            in3 => \N__3514\,
            lcout => \pc.G_12_i_a3_2_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_RNO_0_0_LC_4_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000001010101"
        )
    port map (
            in0 => \N__3515\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__5188\,
            lcout => OPEN,
            ltout => \seq.counter.T8_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_0_LC_4_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1011",
            LUT_INIT => "0001000000000000"
        )
    port map (
            in0 => \N__8551\,
            in1 => \N__4690\,
            in2 => \N__3572\,
            in3 => \N__5366\,
            lcout => \seq_T_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVseq.counter.T_0C_net\,
            ce => 'H',
            sr => \N__7296\
        );

    \pc.program_counter_RNO_2_3_LC_4_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110000000"
        )
    port map (
            in0 => \N__3662\,
            in1 => \N__8548\,
            in2 => \N__3569\,
            in3 => \N__4010\,
            lcout => \pc.N_188_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_1_LC_4_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__3516\,
            lcout => inc,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVseq.counter.T_0C_net\,
            ce => 'H',
            sr => \N__7296\
        );

    \pc.program_counter_RNO_3_3_LC_4_10_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101010100010001"
        )
    port map (
            in0 => \N__8550\,
            in1 => \N__4579\,
            in2 => \_gnd_net_\,
            in3 => \N__4206\,
            lcout => \pc.un1_inc_0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_1_2_LC_4_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100011100000011"
        )
    port map (
            in0 => \N__5760\,
            in1 => \N__5679\,
            in2 => \N__3740\,
            in3 => \N__3820\,
            lcout => OPEN,
            ltout => \pc.G_10_0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_2_LC_4_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101010"
        )
    port map (
            in0 => \N__4088\,
            in1 => \N__3773\,
            in2 => \N__3752\,
            in3 => \N__3749\,
            lcout => \pc.program_counterZ0Z_2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4786\,
            ce => 'H',
            sr => \N__7300\
        );

    \pc.program_counter_RNO_5_2_LC_4_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0101101010101111"
        )
    port map (
            in0 => \N__6162\,
            in1 => \_gnd_net_\,
            in2 => \N__8258\,
            in3 => \N__5990\,
            lcout => \pc.G_10_0_5_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.g0_3_LC_4_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001100110"
        )
    port map (
            in0 => \N__5991\,
            in1 => \N__8257\,
            in2 => \_gnd_net_\,
            in3 => \N__6163\,
            lcout => \ALU_main_N_43_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.un1_A_axb_2_l_ofx_LC_4_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__5992\,
            in1 => \N__8253\,
            in2 => \_gnd_net_\,
            in3 => \N__6161\,
            lcout => \ALU_main.un1_A_axb_2_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_4_2_LC_4_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0110011011001100"
        )
    port map (
            in0 => \N__4833\,
            in1 => \N__3700\,
            in2 => \_gnd_net_\,
            in3 => \N__3666\,
            lcout => \pc.N_10_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.un1_A_cry_0_c_THRU_CRY_0_LC_4_12_0\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__3622\,
            in2 => \N__3626\,
            in3 => \_gnd_net_\,
            lcout => OPEN,
            ltout => OPEN,
            carryin => \bfn_4_12_0_\,
            carryout => \ALU_main.un1_A_cry_0_c_THRU_CO\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.un1_A_cry_0_s_LC_4_12_1\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6060\,
            in2 => \N__4928\,
            in3 => \N__3608\,
            lcout => \un1_A_cry_0_s\,
            ltout => OPEN,
            carryin => \ALU_main.un1_A_cry_0_c_THRU_CO\,
            carryout => \ALU_main.un1_A_cry_0\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.un1_A_cry_0_c_RNIPCLO2_LC_4_12_2\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__6028\,
            in2 => \N__5060\,
            in3 => \N__3605\,
            lcout => \un1_A_cry_0_c_RNIPCLO2\,
            ltout => OPEN,
            carryin => \ALU_main.un1_A_cry_0\,
            carryout => \ALU_main.un1_A_cry_1\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.un1_A_cry_1_c_RNITKPO2_LC_4_12_3\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5989\,
            in2 => \N__3833\,
            in3 => \N__3809\,
            lcout => \un1_A_cry_1_c_RNITKPO2\,
            ltout => OPEN,
            carryin => \ALU_main.un1_A_cry_1\,
            carryout => \ALU_main.un1_A_cry_2\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.un1_A_cry_2_c_RNI1TTO2_LC_4_12_4\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__4919\,
            in2 => \N__5828\,
            in3 => \N__3806\,
            lcout => \un1_A_cry_2_c_RNI1TTO2\,
            ltout => OPEN,
            carryin => \ALU_main.un1_A_cry_2\,
            carryout => \ALU_main.un1_A_cry_3\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.un1_A_cry_3_c_RNI552P2_LC_4_12_5\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5051\,
            in2 => \N__7908\,
            in3 => \N__3803\,
            lcout => \ALU_main.un1_A_cry_3_c_RNI552PZ0Z2\,
            ltout => OPEN,
            carryin => \ALU_main.un1_A_cry_3\,
            carryout => \ALU_main.un1_A_cry_4\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.un1_A_cry_4_c_RNI9D6P2_LC_4_12_6\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5228\,
            in2 => \N__5855\,
            in3 => \N__3800\,
            lcout => \ALU_main.un1_A_cry_4_c_RNI9D6PZ0Z2\,
            ltout => OPEN,
            carryin => \ALU_main.un1_A_cry_4\,
            carryout => \ALU_main.un1_A_cry_5\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.un1_A_cry_5_c_RNIDLAP2_LC_4_12_7\ : LogicCell40
    generic map (
            C_ON => '1',
            SEQ_MODE => "0000",
            LUT_INIT => "1100001100111100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5885\,
            in2 => \N__5912\,
            in3 => \N__3797\,
            lcout => \ALU_main.un1_A_cry_5_c_RNIDLAPZ0Z2\,
            ltout => OPEN,
            carryin => \ALU_main.un1_A_cry_5\,
            carryout => \ALU_main.un1_A_cry_6\,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.un1_A_cry_6_c_RNIP89E2_LC_4_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001011001101001"
        )
    port map (
            in0 => \N__6167\,
            in1 => \N__5866\,
            in2 => \N__6268\,
            in3 => \N__3794\,
            lcout => \ALU_main.un1_A_cry_6_c_RNIP89EZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mem.data_2_7_0__g0_1_LC_4_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__4118\,
            in1 => \N__5748\,
            in2 => \N__4079\,
            in3 => \N__5675\,
            lcout => alu_out_m_1_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.un1_A_cry_5_c_RNI209N9_LC_4_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__5747\,
            in1 => \N__3779\,
            in2 => \N__5924\,
            in3 => \N__5674\,
            lcout => alu_out_m_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.g0_LC_4_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001100110"
        )
    port map (
            in0 => \N__5820\,
            in1 => \N__7833\,
            in2 => \_gnd_net_\,
            in3 => \N__6166\,
            lcout => OPEN,
            ltout => \ALU_main_N_44_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mem.data_2_7_0__g0_0_LC_4_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__5746\,
            in1 => \N__5673\,
            in2 => \N__4121\,
            in3 => \N__4117\,
            lcout => alu_out_m_0_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_0_2_LC_4_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101100010001000"
        )
    port map (
            in0 => \N__8621\,
            in1 => \N__4109\,
            in2 => \N__8434\,
            in3 => \N__4100\,
            lcout => \pc.G_10_0_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.g0_0_LC_4_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001100110"
        )
    port map (
            in0 => \N__5821\,
            in1 => \N__7834\,
            in2 => \_gnd_net_\,
            in3 => \N__6168\,
            lcout => \ALU_main_N_44_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.tbuf.g0_0_1_LC_4_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011001111111111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5823\,
            in2 => \_gnd_net_\,
            in3 => \N__7412\,
            lcout => \pc.tbuf.g0_0_1_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_1_3_LC_4_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100010000000"
        )
    port map (
            in0 => \N__4070\,
            in1 => \N__4061\,
            in2 => \N__4049\,
            in3 => \N__6527\,
            lcout => OPEN,
            ltout => \pc.g0_sn_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_3_LC_4_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111101011001010"
        )
    port map (
            in0 => \N__4031\,
            in1 => \N__3839\,
            in2 => \N__4019\,
            in3 => \N__4016\,
            lcout => \pc.program_counterZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4796\,
            ce => 'H',
            sr => \N__7310\
        );

    \AR.ff4.q_RNILN0E1_LC_4_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000010000000"
        )
    port map (
            in0 => \N__3989\,
            in1 => \N__3971\,
            in2 => \N__3925\,
            in3 => \N__5312\,
            lcout => OPEN,
            ltout => \AR_out_m_3_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.tbuf.g0_0_LC_4_14_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111111011"
        )
    port map (
            in0 => \N__3889\,
            in1 => \N__3848\,
            in2 => \N__3842\,
            in3 => \N__4493\,
            lcout => \pc.g0_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \IR.ff6.q_0_ner_RNIVL0RI_LC_4_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8673\,
            in1 => \N__6079\,
            in2 => \_gnd_net_\,
            in3 => \N__4418\,
            lcout => \N_2_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \IR.ff8.q_0_ner_RNIND22I_LC_4_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110110001000"
        )
    port map (
            in0 => \N__8677\,
            in1 => \N__4388\,
            in2 => \_gnd_net_\,
            in3 => \N__5309\,
            lcout => OPEN,
            ltout => \N_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.q_ret_1_LC_4_15_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0010000000000000"
        )
    port map (
            in0 => \N__5510\,
            in1 => \N__4358\,
            in2 => \N__4340\,
            in3 => \N__4322\,
            lcout => \seq_un1_HLT_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVseq.q_ret_1C_net\,
            ce => 'H',
            sr => \N__7314\
        );

    \seq.counter.T_RNI1G50J_1_LC_4_15_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8674\,
            in2 => \_gnd_net_\,
            in3 => \N__4308\,
            lcout => \seq.un1_HLT_1_reti\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.q_ret_LC_4_16_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "0000000011001100"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8675\,
            in2 => \_gnd_net_\,
            in3 => \N__4309\,
            lcout => \seq.un1_HLT_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVseq.q_retC_net\,
            ce => 'H',
            sr => \N__7319\
        );

    \pc.tbuf.g0_6_LC_5_9_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__8166\,
            in1 => \N__8210\,
            in2 => \N__8129\,
            in3 => \N__8060\,
            lcout => OPEN,
            ltout => \bus_1_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \AR.ff2.q_LC_5_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110001010101010"
        )
    port map (
            in0 => \N__4135\,
            in1 => \N__4692\,
            in2 => \N__4277\,
            in3 => \N__4274\,
            lcout => \AR_out_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVAR.ff2.qC_net\,
            ce => 'H',
            sr => \N__7293\
        );

    \pc.tbuf.out_1_1_iv_0_LC_5_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110101011000000"
        )
    port map (
            in0 => \N__6024\,
            in1 => \N__4214\,
            in2 => \N__4136\,
            in3 => \N__7476\,
            lcout => \pc.tbuf.out_1_1_ivZ0Z_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_3_LC_5_9_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111100000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__4693\,
            lcout => \seq.counter.TZ0Z_3\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVAR.ff2.qC_net\,
            ce => 'H',
            sr => \N__7293\
        );

    \seq.counter.T_RNIPO8O2_3_LC_5_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001001101011111"
        )
    port map (
            in0 => \N__4982\,
            in1 => \N__5096\,
            in2 => \N__5202\,
            in3 => \N__5364\,
            lcout => OPEN,
            ltout => \seq.counter.ACC_LD_0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_RNIIRQM5_4_LC_5_9_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000111111111111"
        )
    port map (
            in0 => \N__5365\,
            in1 => \N__4904\,
            in2 => \N__4874\,
            in3 => \N__6193\,
            lcout => \seq_ACC_LD_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mem.data_2_7_0__g0_i_LC_5_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111101111001111"
        )
    port map (
            in0 => \N__7167\,
            in1 => \N__7108\,
            in2 => \N__7053\,
            in3 => \N__6968\,
            lcout => OPEN,
            ltout => \mem_data_2_7_0__N_11_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.tbuf.g0_7_LC_5_10_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__4871\,
            in1 => \N__4862\,
            in2 => \N__4856\,
            in3 => \N__6537\,
            lcout => \pc.g0_1_0\,
            ltout => \pc.g0_1_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_1_LC_5_10_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011100010"
        )
    port map (
            in0 => \N__4853\,
            in1 => \N__4847\,
            in2 => \N__4841\,
            in3 => \N__8045\,
            lcout => \pc.program_counterZ0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \N__4787\,
            ce => 'H',
            sr => \N__7301\
        );

    \seq.counter.T_0_RNILSL08_0_2_LC_5_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100010000000000"
        )
    port map (
            in0 => \N__4691\,
            in1 => \N__4588\,
            in2 => \N__4430\,
            in3 => \N__4501\,
            lcout => \IR_OE_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.g2_LC_5_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__4980\,
            in1 => \N__5155\,
            in2 => \_gnd_net_\,
            in3 => \N__5014\,
            lcout => \seq.gZ0Z2\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.g0_2_LC_5_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101000100"
        )
    port map (
            in0 => \N__6157\,
            in1 => \N__6014\,
            in2 => \_gnd_net_\,
            in3 => \N__6854\,
            lcout => OPEN,
            ltout => \ALU_main_N_42_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_RNI439M9_4_LC_5_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__5762\,
            in1 => \N__5682\,
            in2 => \N__5045\,
            in3 => \N__5042\,
            lcout => alu_out_m_0_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.g0_1_LC_5_11_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101000100"
        )
    port map (
            in0 => \N__6158\,
            in1 => \N__6050\,
            in2 => \_gnd_net_\,
            in3 => \N__6244\,
            lcout => OPEN,
            ltout => \ALU_main_N_41_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_RNIP3LPB_4_LC_5_11_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010000110000"
        )
    port map (
            in0 => \N__5763\,
            in1 => \N__5683\,
            in2 => \N__5036\,
            in3 => \N__5029\,
            lcout => alu_out_m_0_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.g2_1_LC_5_11_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000010001"
        )
    port map (
            in0 => \N__5015\,
            in1 => \N__4981\,
            in2 => \_gnd_net_\,
            in3 => \N__5156\,
            lcout => \seq.g2Z0Z_1\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.un1_A_axb_0_l_ofx_LC_5_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__6243\,
            in1 => \N__6051\,
            in2 => \_gnd_net_\,
            in3 => \N__6156\,
            lcout => \ALU_main.un1_A_axb_0_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acc.ff6.q_RNI207H1_LC_5_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101000000000"
        )
    port map (
            in0 => \N__5853\,
            in1 => \_gnd_net_\,
            in2 => \_gnd_net_\,
            in3 => \N__7454\,
            lcout => acc_out_m_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.un1_A_axb_3_l_ofx_LC_5_12_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__5822\,
            in1 => \N__7835\,
            in2 => \_gnd_net_\,
            in3 => \N__6164\,
            lcout => \ALU_main.un1_A_axb_3_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.ALU_Out_0_5_LC_5_12_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101000100"
        )
    port map (
            in0 => \N__6165\,
            in1 => \N__5852\,
            in2 => \_gnd_net_\,
            in3 => \N__6359\,
            lcout => OPEN,
            ltout => \ALU_main.N_46_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.un1_A_cry_4_c_RNISJ2N9_LC_5_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0100010011110000"
        )
    port map (
            in0 => \N__5768\,
            in1 => \N__4913\,
            in2 => \N__4907\,
            in3 => \N__5680\,
            lcout => alu_out_m_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.g0_i_a3_0_2_LC_5_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001000000000"
        )
    port map (
            in0 => \N__5504\,
            in1 => \N__5456\,
            in2 => \_gnd_net_\,
            in3 => \N__5406\,
            lcout => OPEN,
            ltout => \seq.g0_i_a3_0Z0Z_2_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_RNI51KH1_4_LC_5_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1101110111011111"
        )
    port map (
            in0 => \N__5363\,
            in1 => \N__5310\,
            in2 => \N__5246\,
            in3 => \N__5243\,
            lcout => \seq_S0_0\,
            ltout => \seq_S0_0_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.un1_A_axb_5_l_ofx_LC_5_12_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5854\,
            in2 => \N__5231\,
            in3 => \N__6358\,
            lcout => \ALU_main.un1_A_axb_5_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \seq.counter.T_RNIR83I4_3_LC_5_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101010001010"
        )
    port map (
            in0 => \N__5203\,
            in1 => \N__5154\,
            in2 => \N__5108\,
            in3 => \N__5092\,
            lcout => \seq_B_LD_0_i\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.un1_A_axb_1_l_ofx_LC_5_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__6029\,
            in1 => \N__6847\,
            in2 => \_gnd_net_\,
            in3 => \N__6159\,
            lcout => \ALU_main.un1_A_axb_1_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_reg.ff5.q_LC_5_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__7951\,
            in1 => \N__7994\,
            in2 => \N__7914\,
            in3 => \N__7456\,
            lcout => b_reg_out_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVb_reg.ff5.qC_net\,
            ce => \N__7781\,
            sr => \N__7311\
        );

    \ALU_main.un1_A_axb_4_l_ofx_LC_5_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1010101001010101"
        )
    port map (
            in0 => \N__6160\,
            in1 => \N__7903\,
            in2 => \_gnd_net_\,
            in3 => \N__6205\,
            lcout => \ALU_main.un1_A_axb_4_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acc.ff7.q_RNI328H1_LC_5_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__5908\,
            in2 => \_gnd_net_\,
            in3 => \N__7455\,
            lcout => acc_out_m_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acc.ff7.q_LC_5_14_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__6821\,
            in1 => \N__6778\,
            in2 => \N__6735\,
            in3 => \N__6535\,
            lcout => acc_out_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacc.ff7.qC_net\,
            ce => \N__5948\,
            sr => \N__7315\
        );

    \ALU_main.ALU_Out_0_6_LC_5_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1001100101000100"
        )
    port map (
            in0 => \N__6191\,
            in1 => \N__5906\,
            in2 => \_gnd_net_\,
            in3 => \N__6704\,
            lcout => \ALU_main.N_47\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.un1_A_axb_6_l_ofx_LC_5_14_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1100110000110011"
        )
    port map (
            in0 => \N__5907\,
            in1 => \N__6703\,
            in2 => \_gnd_net_\,
            in3 => \N__6190\,
            lcout => \ALU_main.un1_A_axb_6_l_ofxZ0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \acc.ff8.q_LC_5_14_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001101"
        )
    port map (
            in0 => \N__6536\,
            in1 => \N__6350\,
            in2 => \N__6891\,
            in3 => \N__6310\,
            lcout => acc_out_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacc.ff7.qC_net\,
            ce => \N__5948\,
            sr => \N__7315\
        );

    \acc.ff6.q_LC_5_14_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__6636\,
            in1 => \N__6683\,
            in2 => \N__6599\,
            in3 => \N__6534\,
            lcout => acc_out_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacc.ff7.qC_net\,
            ce => \N__5948\,
            sr => \N__7315\
        );

    \acc.ff4.q_LC_5_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__7741\,
            in1 => \N__7680\,
            in2 => \N__7619\,
            in3 => \N__7524\,
            lcout => acc_out_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacc.ff7.qC_net\,
            ce => \N__5948\,
            sr => \N__7315\
        );

    \ALU_main.un1_A_cry_3_c_RNIM7SM9_LC_5_15_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0010001011110000"
        )
    port map (
            in0 => \N__5777\,
            in1 => \N__5767\,
            in2 => \N__6095\,
            in3 => \N__5681\,
            lcout => alu_out_m_4,
            ltout => \alu_out_m_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf1.out_1_2_iv_LC_5_15_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111111011111100"
        )
    port map (
            in0 => \N__7910\,
            in1 => \N__7959\,
            in2 => \N__5597\,
            in3 => \N__7457\,
            lcout => bus_4,
            ltout => \bus_4_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \IR.ff5.q_0_ner_RNINVSHI_LC_5_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111001111000000"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \N__8676\,
            in2 => \N__5567\,
            in3 => \N__5563\,
            lcout => \N_4_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \ALU_main.ALU_Out_0_4_LC_5_15_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1000100001100110"
        )
    port map (
            in0 => \N__7909\,
            in1 => \N__6209\,
            in2 => \_gnd_net_\,
            in3 => \N__6192\,
            lcout => \ALU_main.N_45\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \buf1.out_1_1_iv_LC_5_15_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "1111101011111011"
        )
    port map (
            in0 => \N__6635\,
            in1 => \N__6600\,
            in2 => \N__6690\,
            in3 => \N__6551\,
            lcout => bus_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \IR.ff2.q_ner_LC_6_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__8211\,
            in1 => \N__8168\,
            in2 => \N__8121\,
            in3 => \N__8064\,
            lcout => ir_out_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVIR.ff2.q_nerC_net\,
            ce => \N__8678\,
            sr => \N__7297\
        );

    \IR.ff3.q_ner_LC_6_9_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__8425\,
            in1 => \N__8457\,
            in2 => \N__8368\,
            in3 => \N__8293\,
            lcout => ir_out_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVIR.ff2.q_nerC_net\,
            ce => \N__8678\,
            sr => \N__7297\
        );

    \acc.ff1.q_LC_6_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__8919\,
            in1 => \N__8731\,
            in2 => \N__8860\,
            in3 => \N__8794\,
            lcout => acc_out_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacc.ff1.qC_net\,
            ce => \N__5947\,
            sr => \N__7305\
        );

    \acc.ff2.q_LC_6_10_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__8167\,
            in1 => \N__8229\,
            in2 => \N__8122\,
            in3 => \N__8053\,
            lcout => acc_out_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacc.ff1.qC_net\,
            ce => \N__5947\,
            sr => \N__7305\
        );

    \acc.ff3.q_LC_6_10_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__8306\,
            in1 => \N__8411\,
            in2 => \N__8373\,
            in3 => \N__8478\,
            lcout => acc_out_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacc.ff1.qC_net\,
            ce => \N__5947\,
            sr => \N__7305\
        );

    \acc.ff5.q_LC_6_10_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__8003\,
            in1 => \N__7960\,
            in2 => \N__7904\,
            in3 => \N__7479\,
            lcout => acc_out_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVacc.ff1.qC_net\,
            ce => \N__5947\,
            sr => \N__7305\
        );

    \mar.ff4.q_ner_LC_6_11_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__7748\,
            in1 => \N__7678\,
            in2 => \N__7630\,
            in3 => \N__7546\,
            lcout => mar_out_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVmar.ff4.q_nerC_net\,
            ce => \N__6383\,
            sr => \N__7308\
        );

    \mar.ff3.q_ner_LC_6_11_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__8426\,
            in1 => \N__8307\,
            in2 => \N__8374\,
            in3 => \N__8479\,
            lcout => mar_out_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVmar.ff4.q_nerC_net\,
            ce => \N__6383\,
            sr => \N__7308\
        );

    \mar.ff2.q_ner_LC_6_11_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__8236\,
            in1 => \N__8169\,
            in2 => \N__8130\,
            in3 => \N__8052\,
            lcout => mar_out_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVmar.ff4.q_nerC_net\,
            ce => \N__6383\,
            sr => \N__7308\
        );

    \b_reg.ff6.q_LC_6_12_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__6670\,
            in1 => \N__6634\,
            in2 => \N__6598\,
            in3 => \N__6555\,
            lcout => b_reg_out_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVb_reg.ff6.qC_net\,
            ce => \N__7804\,
            sr => \N__7312\
        );

    \b_reg.ff8.q_LC_6_12_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001101"
        )
    port map (
            in0 => \N__6556\,
            in1 => \N__6346\,
            in2 => \N__6890\,
            in3 => \N__6311\,
            lcout => b_reg_out_7,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVb_reg.ff6.qC_net\,
            ce => \N__7804\,
            sr => \N__7312\
        );

    \b_reg.ff1.q_LC_6_12_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__8927\,
            in1 => \N__8848\,
            in2 => \N__8755\,
            in3 => \N__8795\,
            lcout => b_reg_out_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVb_reg.ff6.qC_net\,
            ce => \N__7804\,
            sr => \N__7312\
        );

    \mem.data_2_7_0__m18_LC_6_13_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111000101111"
        )
    port map (
            in0 => \N__6962\,
            in1 => \N__7176\,
            in2 => \N__7128\,
            in3 => \N__7029\,
            lcout => OPEN,
            ltout => \mem.i2_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mem.data_2_7_0__i2_mux_i_m_LC_6_13_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0000000000001111"
        )
    port map (
            in0 => \_gnd_net_\,
            in1 => \_gnd_net_\,
            in2 => \N__6224\,
            in3 => \N__6553\,
            lcout => \mem_data_2_7_0__i2_mux_i_m\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \pc.program_counter_RNO_10_0_LC_6_13_3\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111111110011011"
        )
    port map (
            in0 => \N__7175\,
            in1 => \N__7109\,
            in2 => \N__7045\,
            in3 => \N__6960\,
            lcout => \pc.N_7\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mem.data_2_7_0__m20_LC_6_13_4\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0011111111010111"
        )
    port map (
            in0 => \N__6961\,
            in1 => \N__7177\,
            in2 => \N__7127\,
            in3 => \N__7028\,
            lcout => m20,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \mem.data_2_7_0__m22_LC_6_13_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0111010101110111"
        )
    port map (
            in0 => \N__7178\,
            in1 => \N__7114\,
            in2 => \N__7046\,
            in3 => \N__6963\,
            lcout => \mem_data_2_7_0__N_29_mux\,
            ltout => \mem_data_2_7_0__N_29_mux_cascade_\,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \out_reg.ff7.q_LC_6_13_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001101"
        )
    port map (
            in0 => \N__6554\,
            in1 => \N__6820\,
            in2 => \N__7208\,
            in3 => \N__6782\,
            lcout => out_c_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVout_reg.ff7.qC_net\,
            ce => \N__7473\,
            sr => \N__7316\
        );

    \mem.data_2_7_0__m26_LC_6_13_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "0000",
            LUT_INIT => "0001111011111001"
        )
    port map (
            in0 => \N__7179\,
            in1 => \N__7113\,
            in2 => \N__7047\,
            in3 => \N__6964\,
            lcout => \mem_data_2_7_0__i2_mux_0\,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \_gnd_net_\,
            ce => 'H',
            sr => \_gnd_net_\
        );

    \b_reg.ff2.q_LC_6_14_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__8237\,
            in1 => \N__8183\,
            in2 => \N__8138\,
            in3 => \N__8065\,
            lcout => b_reg_out_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVb_reg.ff2.qC_net\,
            ce => \N__7811\,
            sr => \N__7320\
        );

    \b_reg.ff7.q_LC_6_14_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__6822\,
            in1 => \N__6790\,
            in2 => \N__6734\,
            in3 => \N__6557\,
            lcout => b_reg_out_6,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVb_reg.ff2.qC_net\,
            ce => \N__7811\,
            sr => \N__7320\
        );

    \out_reg.ff6.q_LC_6_15_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1110111011101111"
        )
    port map (
            in0 => \N__6691\,
            in1 => \N__6637\,
            in2 => \N__6604\,
            in3 => \N__6552\,
            lcout => out_c_5,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVout_reg.ff6.qC_net\,
            ce => \N__7474\,
            sr => \N__7322\
        );

    \out_reg.ff3.q_LC_7_9_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111001110"
        )
    port map (
            in0 => \N__8412\,
            in1 => \N__8468\,
            in2 => \N__8369\,
            in3 => \N__8309\,
            lcout => out_c_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVout_reg.ff3.qC_net\,
            ce => \N__7484\,
            sr => \N__7302\
        );

    \out_reg.ff1.q_LC_7_9_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__8909\,
            in1 => \N__8732\,
            in2 => \N__8879\,
            in3 => \N__8816\,
            lcout => out_c_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVout_reg.ff3.qC_net\,
            ce => \N__7484\,
            sr => \N__7302\
        );

    \IR.ff1.q_ner_LC_7_10_0\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110111010"
        )
    port map (
            in0 => \N__8926\,
            in1 => \N__8873\,
            in2 => \N__8748\,
            in3 => \N__8815\,
            lcout => ir_out_0,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVIR.ff1.q_nerC_net\,
            ce => \N__8679\,
            sr => \N__7309\
        );

    \b_reg.ff3.q_LC_7_11_1\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111110101110"
        )
    port map (
            in0 => \N__8480\,
            in1 => \N__8427\,
            in2 => \N__8375\,
            in3 => \N__8308\,
            lcout => b_reg_out_2,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVb_reg.ff3.qC_net\,
            ce => \N__7803\,
            sr => \N__7313\
        );

    \out_reg.ff2.q_LC_7_12_5\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111011100"
        )
    port map (
            in0 => \N__8228\,
            in1 => \N__8182\,
            in2 => \N__8137\,
            in3 => \N__8066\,
            lcout => out_c_1,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVout_reg.ff2.qC_net\,
            ce => \N__7478\,
            sr => \N__7317\
        );

    \out_reg.ff5.q_LC_7_12_6\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111011101110"
        )
    port map (
            in0 => \N__8002\,
            in1 => \N__7952\,
            in2 => \N__7915\,
            in3 => \N__7477\,
            lcout => out_c_4,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVout_reg.ff2.qC_net\,
            ce => \N__7478\,
            sr => \N__7317\
        );

    \b_reg.ff4.q_LC_7_13_2\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__7750\,
            in1 => \N__7685\,
            in2 => \N__7620\,
            in3 => \N__7540\,
            lcout => b_reg_out_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVb_reg.ff4.qC_net\,
            ce => \N__7793\,
            sr => \N__7321\
        );

    \out_reg.ff4.q_LC_8_11_7\ : LogicCell40
    generic map (
            C_ON => '0',
            SEQ_MODE => "1010",
            LUT_INIT => "1111111111101111"
        )
    port map (
            in0 => \N__7754\,
            in1 => \N__7679\,
            in2 => \N__7631\,
            in3 => \N__7547\,
            lcout => out_c_3,
            ltout => OPEN,
            carryin => \_gnd_net_\,
            carryout => OPEN,
            clk => \INVout_reg.ff4.qC_net\,
            ce => \N__7475\,
            sr => \N__7318\
        );
end \INTERFACE\;
