// ******************************************************************************

// iCEcube Netlister

// Version:            2020.12.27943

// Build Date:         Dec  9 2020 18:18:12

// File Generated:     Dec 13 2023 19:34:34

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "test" view "INTERFACE"

module test (
    LED4,
    LED2,
    LED5,
    LED3,
    LED1);

    output LED4;
    output LED2;
    output LED5;
    output LED3;
    output LED1;

    wire N__9920;
    wire N__9919;
    wire N__9918;
    wire N__9911;
    wire N__9910;
    wire N__9909;
    wire N__9902;
    wire N__9901;
    wire N__9900;
    wire N__9893;
    wire N__9892;
    wire N__9891;
    wire N__9884;
    wire N__9883;
    wire N__9882;
    wire N__9865;
    wire N__9862;
    wire N__9859;
    wire N__9856;
    wire N__9853;
    wire N__9852;
    wire N__9851;
    wire N__9850;
    wire N__9847;
    wire N__9844;
    wire N__9841;
    wire N__9840;
    wire N__9837;
    wire N__9836;
    wire N__9829;
    wire N__9826;
    wire N__9823;
    wire N__9820;
    wire N__9815;
    wire N__9808;
    wire N__9805;
    wire N__9804;
    wire N__9803;
    wire N__9802;
    wire N__9799;
    wire N__9796;
    wire N__9793;
    wire N__9790;
    wire N__9785;
    wire N__9782;
    wire N__9779;
    wire N__9772;
    wire N__9771;
    wire N__9768;
    wire N__9767;
    wire N__9764;
    wire N__9763;
    wire N__9760;
    wire N__9757;
    wire N__9754;
    wire N__9751;
    wire N__9748;
    wire N__9743;
    wire N__9740;
    wire N__9739;
    wire N__9736;
    wire N__9733;
    wire N__9730;
    wire N__9727;
    wire N__9718;
    wire N__9715;
    wire N__9714;
    wire N__9713;
    wire N__9712;
    wire N__9711;
    wire N__9708;
    wire N__9705;
    wire N__9702;
    wire N__9697;
    wire N__9692;
    wire N__9687;
    wire N__9684;
    wire N__9681;
    wire N__9676;
    wire N__9675;
    wire N__9672;
    wire N__9671;
    wire N__9670;
    wire N__9667;
    wire N__9666;
    wire N__9665;
    wire N__9656;
    wire N__9655;
    wire N__9654;
    wire N__9653;
    wire N__9652;
    wire N__9651;
    wire N__9650;
    wire N__9645;
    wire N__9642;
    wire N__9637;
    wire N__9632;
    wire N__9629;
    wire N__9626;
    wire N__9613;
    wire N__9612;
    wire N__9611;
    wire N__9610;
    wire N__9609;
    wire N__9608;
    wire N__9607;
    wire N__9604;
    wire N__9601;
    wire N__9600;
    wire N__9597;
    wire N__9594;
    wire N__9591;
    wire N__9590;
    wire N__9589;
    wire N__9586;
    wire N__9577;
    wire N__9572;
    wire N__9571;
    wire N__9566;
    wire N__9561;
    wire N__9556;
    wire N__9553;
    wire N__9544;
    wire N__9543;
    wire N__9540;
    wire N__9539;
    wire N__9536;
    wire N__9535;
    wire N__9530;
    wire N__9527;
    wire N__9526;
    wire N__9525;
    wire N__9524;
    wire N__9523;
    wire N__9522;
    wire N__9521;
    wire N__9520;
    wire N__9517;
    wire N__9512;
    wire N__9509;
    wire N__9500;
    wire N__9495;
    wire N__9490;
    wire N__9481;
    wire N__9478;
    wire N__9475;
    wire N__9472;
    wire N__9469;
    wire N__9468;
    wire N__9465;
    wire N__9464;
    wire N__9461;
    wire N__9460;
    wire N__9459;
    wire N__9458;
    wire N__9455;
    wire N__9452;
    wire N__9449;
    wire N__9446;
    wire N__9441;
    wire N__9436;
    wire N__9427;
    wire N__9424;
    wire N__9421;
    wire N__9420;
    wire N__9419;
    wire N__9416;
    wire N__9413;
    wire N__9410;
    wire N__9403;
    wire N__9402;
    wire N__9401;
    wire N__9400;
    wire N__9397;
    wire N__9396;
    wire N__9395;
    wire N__9394;
    wire N__9393;
    wire N__9390;
    wire N__9387;
    wire N__9384;
    wire N__9381;
    wire N__9378;
    wire N__9373;
    wire N__9370;
    wire N__9367;
    wire N__9364;
    wire N__9363;
    wire N__9362;
    wire N__9357;
    wire N__9356;
    wire N__9353;
    wire N__9350;
    wire N__9345;
    wire N__9342;
    wire N__9337;
    wire N__9334;
    wire N__9331;
    wire N__9324;
    wire N__9313;
    wire N__9310;
    wire N__9309;
    wire N__9306;
    wire N__9303;
    wire N__9298;
    wire N__9297;
    wire N__9294;
    wire N__9291;
    wire N__9286;
    wire N__9283;
    wire N__9280;
    wire N__9279;
    wire N__9278;
    wire N__9275;
    wire N__9270;
    wire N__9265;
    wire N__9262;
    wire N__9259;
    wire N__9258;
    wire N__9255;
    wire N__9252;
    wire N__9247;
    wire N__9244;
    wire N__9241;
    wire N__9240;
    wire N__9239;
    wire N__9236;
    wire N__9233;
    wire N__9230;
    wire N__9227;
    wire N__9224;
    wire N__9221;
    wire N__9220;
    wire N__9217;
    wire N__9212;
    wire N__9209;
    wire N__9206;
    wire N__9201;
    wire N__9196;
    wire N__9195;
    wire N__9194;
    wire N__9191;
    wire N__9188;
    wire N__9185;
    wire N__9182;
    wire N__9179;
    wire N__9176;
    wire N__9175;
    wire N__9172;
    wire N__9169;
    wire N__9166;
    wire N__9163;
    wire N__9158;
    wire N__9155;
    wire N__9152;
    wire N__9147;
    wire N__9144;
    wire N__9139;
    wire N__9138;
    wire N__9137;
    wire N__9134;
    wire N__9133;
    wire N__9130;
    wire N__9127;
    wire N__9124;
    wire N__9123;
    wire N__9120;
    wire N__9117;
    wire N__9114;
    wire N__9111;
    wire N__9110;
    wire N__9107;
    wire N__9104;
    wire N__9101;
    wire N__9098;
    wire N__9095;
    wire N__9092;
    wire N__9079;
    wire N__9078;
    wire N__9077;
    wire N__9076;
    wire N__9075;
    wire N__9074;
    wire N__9073;
    wire N__9072;
    wire N__9071;
    wire N__9068;
    wire N__9065;
    wire N__9058;
    wire N__9055;
    wire N__9054;
    wire N__9053;
    wire N__9050;
    wire N__9047;
    wire N__9046;
    wire N__9045;
    wire N__9044;
    wire N__9043;
    wire N__9042;
    wire N__9039;
    wire N__9038;
    wire N__9037;
    wire N__9034;
    wire N__9033;
    wire N__9032;
    wire N__9029;
    wire N__9026;
    wire N__9023;
    wire N__9020;
    wire N__9017;
    wire N__9012;
    wire N__9009;
    wire N__9006;
    wire N__9005;
    wire N__9002;
    wire N__8995;
    wire N__8992;
    wire N__8989;
    wire N__8986;
    wire N__8985;
    wire N__8984;
    wire N__8981;
    wire N__8978;
    wire N__8977;
    wire N__8976;
    wire N__8975;
    wire N__8974;
    wire N__8973;
    wire N__8972;
    wire N__8971;
    wire N__8968;
    wire N__8961;
    wire N__8954;
    wire N__8951;
    wire N__8948;
    wire N__8941;
    wire N__8938;
    wire N__8935;
    wire N__8932;
    wire N__8929;
    wire N__8924;
    wire N__8923;
    wire N__8920;
    wire N__8917;
    wire N__8908;
    wire N__8905;
    wire N__8902;
    wire N__8897;
    wire N__8892;
    wire N__8889;
    wire N__8880;
    wire N__8877;
    wire N__8874;
    wire N__8851;
    wire N__8850;
    wire N__8849;
    wire N__8848;
    wire N__8847;
    wire N__8846;
    wire N__8845;
    wire N__8844;
    wire N__8843;
    wire N__8842;
    wire N__8833;
    wire N__8828;
    wire N__8827;
    wire N__8822;
    wire N__8817;
    wire N__8812;
    wire N__8809;
    wire N__8800;
    wire N__8799;
    wire N__8796;
    wire N__8793;
    wire N__8790;
    wire N__8787;
    wire N__8784;
    wire N__8781;
    wire N__8778;
    wire N__8773;
    wire N__8770;
    wire N__8769;
    wire N__8768;
    wire N__8767;
    wire N__8766;
    wire N__8765;
    wire N__8762;
    wire N__8761;
    wire N__8758;
    wire N__8757;
    wire N__8756;
    wire N__8753;
    wire N__8750;
    wire N__8745;
    wire N__8744;
    wire N__8741;
    wire N__8736;
    wire N__8733;
    wire N__8730;
    wire N__8727;
    wire N__8724;
    wire N__8721;
    wire N__8718;
    wire N__8717;
    wire N__8716;
    wire N__8715;
    wire N__8710;
    wire N__8707;
    wire N__8704;
    wire N__8695;
    wire N__8692;
    wire N__8689;
    wire N__8686;
    wire N__8683;
    wire N__8676;
    wire N__8673;
    wire N__8670;
    wire N__8659;
    wire N__8658;
    wire N__8657;
    wire N__8656;
    wire N__8655;
    wire N__8654;
    wire N__8651;
    wire N__8648;
    wire N__8643;
    wire N__8638;
    wire N__8635;
    wire N__8634;
    wire N__8633;
    wire N__8630;
    wire N__8627;
    wire N__8624;
    wire N__8621;
    wire N__8616;
    wire N__8611;
    wire N__8602;
    wire N__8601;
    wire N__8598;
    wire N__8597;
    wire N__8594;
    wire N__8591;
    wire N__8586;
    wire N__8581;
    wire N__8580;
    wire N__8579;
    wire N__8578;
    wire N__8577;
    wire N__8576;
    wire N__8575;
    wire N__8574;
    wire N__8569;
    wire N__8566;
    wire N__8559;
    wire N__8556;
    wire N__8553;
    wire N__8552;
    wire N__8551;
    wire N__8550;
    wire N__8549;
    wire N__8546;
    wire N__8541;
    wire N__8536;
    wire N__8531;
    wire N__8528;
    wire N__8525;
    wire N__8522;
    wire N__8515;
    wire N__8510;
    wire N__8503;
    wire N__8500;
    wire N__8497;
    wire N__8496;
    wire N__8495;
    wire N__8492;
    wire N__8489;
    wire N__8488;
    wire N__8485;
    wire N__8482;
    wire N__8479;
    wire N__8478;
    wire N__8477;
    wire N__8474;
    wire N__8471;
    wire N__8466;
    wire N__8465;
    wire N__8464;
    wire N__8461;
    wire N__8458;
    wire N__8455;
    wire N__8450;
    wire N__8445;
    wire N__8442;
    wire N__8431;
    wire N__8430;
    wire N__8427;
    wire N__8426;
    wire N__8423;
    wire N__8420;
    wire N__8417;
    wire N__8416;
    wire N__8411;
    wire N__8408;
    wire N__8405;
    wire N__8404;
    wire N__8401;
    wire N__8398;
    wire N__8393;
    wire N__8386;
    wire N__8385;
    wire N__8384;
    wire N__8383;
    wire N__8382;
    wire N__8379;
    wire N__8376;
    wire N__8375;
    wire N__8372;
    wire N__8369;
    wire N__8366;
    wire N__8361;
    wire N__8360;
    wire N__8359;
    wire N__8356;
    wire N__8353;
    wire N__8350;
    wire N__8347;
    wire N__8344;
    wire N__8341;
    wire N__8338;
    wire N__8335;
    wire N__8332;
    wire N__8329;
    wire N__8324;
    wire N__8321;
    wire N__8308;
    wire N__8305;
    wire N__8302;
    wire N__8301;
    wire N__8298;
    wire N__8295;
    wire N__8290;
    wire N__8287;
    wire N__8286;
    wire N__8283;
    wire N__8282;
    wire N__8281;
    wire N__8280;
    wire N__8279;
    wire N__8278;
    wire N__8275;
    wire N__8274;
    wire N__8273;
    wire N__8272;
    wire N__8271;
    wire N__8268;
    wire N__8265;
    wire N__8262;
    wire N__8261;
    wire N__8260;
    wire N__8257;
    wire N__8254;
    wire N__8253;
    wire N__8250;
    wire N__8247;
    wire N__8242;
    wire N__8239;
    wire N__8236;
    wire N__8229;
    wire N__8226;
    wire N__8223;
    wire N__8218;
    wire N__8215;
    wire N__8210;
    wire N__8205;
    wire N__8200;
    wire N__8197;
    wire N__8194;
    wire N__8191;
    wire N__8188;
    wire N__8183;
    wire N__8178;
    wire N__8175;
    wire N__8170;
    wire N__8161;
    wire N__8158;
    wire N__8157;
    wire N__8154;
    wire N__8151;
    wire N__8148;
    wire N__8145;
    wire N__8140;
    wire N__8137;
    wire N__8134;
    wire N__8131;
    wire N__8128;
    wire N__8125;
    wire N__8122;
    wire N__8121;
    wire N__8118;
    wire N__8115;
    wire N__8112;
    wire N__8109;
    wire N__8108;
    wire N__8103;
    wire N__8100;
    wire N__8099;
    wire N__8098;
    wire N__8095;
    wire N__8092;
    wire N__8089;
    wire N__8086;
    wire N__8077;
    wire N__8074;
    wire N__8073;
    wire N__8070;
    wire N__8067;
    wire N__8066;
    wire N__8063;
    wire N__8060;
    wire N__8057;
    wire N__8050;
    wire N__8047;
    wire N__8044;
    wire N__8043;
    wire N__8038;
    wire N__8035;
    wire N__8032;
    wire N__8031;
    wire N__8028;
    wire N__8027;
    wire N__8024;
    wire N__8023;
    wire N__8020;
    wire N__8017;
    wire N__8014;
    wire N__8011;
    wire N__8008;
    wire N__8005;
    wire N__8002;
    wire N__7999;
    wire N__7996;
    wire N__7987;
    wire N__7986;
    wire N__7985;
    wire N__7982;
    wire N__7979;
    wire N__7976;
    wire N__7975;
    wire N__7974;
    wire N__7971;
    wire N__7966;
    wire N__7965;
    wire N__7962;
    wire N__7959;
    wire N__7954;
    wire N__7949;
    wire N__7946;
    wire N__7939;
    wire N__7936;
    wire N__7935;
    wire N__7934;
    wire N__7933;
    wire N__7930;
    wire N__7929;
    wire N__7926;
    wire N__7921;
    wire N__7918;
    wire N__7915;
    wire N__7912;
    wire N__7909;
    wire N__7904;
    wire N__7899;
    wire N__7894;
    wire N__7893;
    wire N__7892;
    wire N__7889;
    wire N__7886;
    wire N__7883;
    wire N__7880;
    wire N__7877;
    wire N__7874;
    wire N__7873;
    wire N__7872;
    wire N__7869;
    wire N__7864;
    wire N__7859;
    wire N__7852;
    wire N__7849;
    wire N__7846;
    wire N__7843;
    wire N__7840;
    wire N__7837;
    wire N__7836;
    wire N__7833;
    wire N__7830;
    wire N__7827;
    wire N__7824;
    wire N__7821;
    wire N__7818;
    wire N__7813;
    wire N__7810;
    wire N__7807;
    wire N__7804;
    wire N__7803;
    wire N__7800;
    wire N__7797;
    wire N__7794;
    wire N__7791;
    wire N__7786;
    wire N__7783;
    wire N__7782;
    wire N__7781;
    wire N__7780;
    wire N__7779;
    wire N__7776;
    wire N__7773;
    wire N__7770;
    wire N__7765;
    wire N__7764;
    wire N__7763;
    wire N__7762;
    wire N__7761;
    wire N__7760;
    wire N__7759;
    wire N__7758;
    wire N__7755;
    wire N__7748;
    wire N__7745;
    wire N__7742;
    wire N__7739;
    wire N__7736;
    wire N__7733;
    wire N__7728;
    wire N__7725;
    wire N__7722;
    wire N__7715;
    wire N__7708;
    wire N__7699;
    wire N__7696;
    wire N__7693;
    wire N__7692;
    wire N__7689;
    wire N__7688;
    wire N__7685;
    wire N__7684;
    wire N__7681;
    wire N__7680;
    wire N__7677;
    wire N__7674;
    wire N__7671;
    wire N__7668;
    wire N__7665;
    wire N__7662;
    wire N__7657;
    wire N__7652;
    wire N__7645;
    wire N__7644;
    wire N__7643;
    wire N__7640;
    wire N__7637;
    wire N__7636;
    wire N__7633;
    wire N__7630;
    wire N__7627;
    wire N__7624;
    wire N__7623;
    wire N__7620;
    wire N__7617;
    wire N__7612;
    wire N__7609;
    wire N__7606;
    wire N__7597;
    wire N__7596;
    wire N__7593;
    wire N__7590;
    wire N__7589;
    wire N__7586;
    wire N__7583;
    wire N__7580;
    wire N__7579;
    wire N__7576;
    wire N__7571;
    wire N__7568;
    wire N__7567;
    wire N__7562;
    wire N__7559;
    wire N__7556;
    wire N__7549;
    wire N__7548;
    wire N__7547;
    wire N__7544;
    wire N__7541;
    wire N__7538;
    wire N__7535;
    wire N__7532;
    wire N__7529;
    wire N__7526;
    wire N__7523;
    wire N__7516;
    wire N__7515;
    wire N__7514;
    wire N__7511;
    wire N__7510;
    wire N__7507;
    wire N__7504;
    wire N__7503;
    wire N__7500;
    wire N__7497;
    wire N__7494;
    wire N__7491;
    wire N__7488;
    wire N__7487;
    wire N__7482;
    wire N__7481;
    wire N__7476;
    wire N__7473;
    wire N__7470;
    wire N__7467;
    wire N__7464;
    wire N__7461;
    wire N__7458;
    wire N__7455;
    wire N__7450;
    wire N__7447;
    wire N__7444;
    wire N__7439;
    wire N__7432;
    wire N__7429;
    wire N__7428;
    wire N__7425;
    wire N__7422;
    wire N__7421;
    wire N__7420;
    wire N__7419;
    wire N__7418;
    wire N__7417;
    wire N__7416;
    wire N__7415;
    wire N__7414;
    wire N__7413;
    wire N__7412;
    wire N__7407;
    wire N__7406;
    wire N__7405;
    wire N__7404;
    wire N__7403;
    wire N__7402;
    wire N__7401;
    wire N__7392;
    wire N__7387;
    wire N__7386;
    wire N__7383;
    wire N__7378;
    wire N__7375;
    wire N__7372;
    wire N__7369;
    wire N__7364;
    wire N__7361;
    wire N__7360;
    wire N__7357;
    wire N__7354;
    wire N__7351;
    wire N__7348;
    wire N__7345;
    wire N__7340;
    wire N__7329;
    wire N__7328;
    wire N__7327;
    wire N__7324;
    wire N__7321;
    wire N__7312;
    wire N__7311;
    wire N__7310;
    wire N__7309;
    wire N__7308;
    wire N__7305;
    wire N__7302;
    wire N__7297;
    wire N__7294;
    wire N__7291;
    wire N__7288;
    wire N__7285;
    wire N__7278;
    wire N__7269;
    wire N__7258;
    wire N__7255;
    wire N__7254;
    wire N__7251;
    wire N__7248;
    wire N__7247;
    wire N__7244;
    wire N__7239;
    wire N__7238;
    wire N__7237;
    wire N__7234;
    wire N__7231;
    wire N__7228;
    wire N__7225;
    wire N__7222;
    wire N__7217;
    wire N__7210;
    wire N__7209;
    wire N__7206;
    wire N__7203;
    wire N__7200;
    wire N__7197;
    wire N__7192;
    wire N__7189;
    wire N__7186;
    wire N__7185;
    wire N__7182;
    wire N__7179;
    wire N__7174;
    wire N__7171;
    wire N__7168;
    wire N__7167;
    wire N__7164;
    wire N__7163;
    wire N__7160;
    wire N__7157;
    wire N__7154;
    wire N__7151;
    wire N__7148;
    wire N__7141;
    wire N__7140;
    wire N__7139;
    wire N__7136;
    wire N__7133;
    wire N__7132;
    wire N__7129;
    wire N__7126;
    wire N__7123;
    wire N__7120;
    wire N__7117;
    wire N__7114;
    wire N__7109;
    wire N__7102;
    wire N__7099;
    wire N__7096;
    wire N__7093;
    wire N__7090;
    wire N__7087;
    wire N__7084;
    wire N__7081;
    wire N__7078;
    wire N__7075;
    wire N__7072;
    wire N__7069;
    wire N__7066;
    wire N__7063;
    wire N__7060;
    wire N__7059;
    wire N__7056;
    wire N__7053;
    wire N__7050;
    wire N__7049;
    wire N__7046;
    wire N__7043;
    wire N__7040;
    wire N__7033;
    wire N__7032;
    wire N__7031;
    wire N__7030;
    wire N__7029;
    wire N__7028;
    wire N__7027;
    wire N__7024;
    wire N__7021;
    wire N__7020;
    wire N__7019;
    wire N__7016;
    wire N__7013;
    wire N__7010;
    wire N__7007;
    wire N__7004;
    wire N__7001;
    wire N__6998;
    wire N__6995;
    wire N__6990;
    wire N__6987;
    wire N__6982;
    wire N__6979;
    wire N__6976;
    wire N__6971;
    wire N__6966;
    wire N__6955;
    wire N__6952;
    wire N__6949;
    wire N__6946;
    wire N__6943;
    wire N__6942;
    wire N__6939;
    wire N__6936;
    wire N__6935;
    wire N__6934;
    wire N__6931;
    wire N__6928;
    wire N__6927;
    wire N__6926;
    wire N__6925;
    wire N__6922;
    wire N__6919;
    wire N__6916;
    wire N__6913;
    wire N__6908;
    wire N__6905;
    wire N__6892;
    wire N__6889;
    wire N__6886;
    wire N__6885;
    wire N__6884;
    wire N__6881;
    wire N__6878;
    wire N__6875;
    wire N__6874;
    wire N__6869;
    wire N__6866;
    wire N__6863;
    wire N__6860;
    wire N__6857;
    wire N__6854;
    wire N__6847;
    wire N__6844;
    wire N__6841;
    wire N__6838;
    wire N__6835;
    wire N__6834;
    wire N__6831;
    wire N__6828;
    wire N__6825;
    wire N__6822;
    wire N__6817;
    wire N__6814;
    wire N__6811;
    wire N__6808;
    wire N__6805;
    wire N__6802;
    wire N__6799;
    wire N__6798;
    wire N__6795;
    wire N__6792;
    wire N__6789;
    wire N__6786;
    wire N__6783;
    wire N__6780;
    wire N__6775;
    wire N__6774;
    wire N__6773;
    wire N__6772;
    wire N__6769;
    wire N__6768;
    wire N__6767;
    wire N__6766;
    wire N__6763;
    wire N__6762;
    wire N__6761;
    wire N__6760;
    wire N__6755;
    wire N__6754;
    wire N__6753;
    wire N__6752;
    wire N__6749;
    wire N__6746;
    wire N__6743;
    wire N__6740;
    wire N__6737;
    wire N__6732;
    wire N__6729;
    wire N__6726;
    wire N__6723;
    wire N__6718;
    wire N__6713;
    wire N__6706;
    wire N__6703;
    wire N__6700;
    wire N__6693;
    wire N__6690;
    wire N__6685;
    wire N__6680;
    wire N__6673;
    wire N__6672;
    wire N__6669;
    wire N__6668;
    wire N__6665;
    wire N__6660;
    wire N__6657;
    wire N__6654;
    wire N__6653;
    wire N__6650;
    wire N__6647;
    wire N__6644;
    wire N__6637;
    wire N__6636;
    wire N__6635;
    wire N__6628;
    wire N__6625;
    wire N__6622;
    wire N__6621;
    wire N__6620;
    wire N__6619;
    wire N__6618;
    wire N__6617;
    wire N__6616;
    wire N__6615;
    wire N__6614;
    wire N__6611;
    wire N__6610;
    wire N__6607;
    wire N__6604;
    wire N__6603;
    wire N__6600;
    wire N__6597;
    wire N__6594;
    wire N__6591;
    wire N__6586;
    wire N__6583;
    wire N__6582;
    wire N__6581;
    wire N__6580;
    wire N__6577;
    wire N__6572;
    wire N__6569;
    wire N__6566;
    wire N__6563;
    wire N__6560;
    wire N__6557;
    wire N__6554;
    wire N__6551;
    wire N__6548;
    wire N__6543;
    wire N__6540;
    wire N__6537;
    wire N__6534;
    wire N__6531;
    wire N__6516;
    wire N__6505;
    wire N__6502;
    wire N__6501;
    wire N__6500;
    wire N__6499;
    wire N__6498;
    wire N__6497;
    wire N__6496;
    wire N__6493;
    wire N__6492;
    wire N__6489;
    wire N__6486;
    wire N__6479;
    wire N__6476;
    wire N__6475;
    wire N__6474;
    wire N__6471;
    wire N__6468;
    wire N__6467;
    wire N__6464;
    wire N__6463;
    wire N__6460;
    wire N__6457;
    wire N__6456;
    wire N__6453;
    wire N__6450;
    wire N__6447;
    wire N__6442;
    wire N__6439;
    wire N__6436;
    wire N__6433;
    wire N__6428;
    wire N__6425;
    wire N__6406;
    wire N__6403;
    wire N__6402;
    wire N__6399;
    wire N__6396;
    wire N__6395;
    wire N__6392;
    wire N__6389;
    wire N__6388;
    wire N__6385;
    wire N__6380;
    wire N__6377;
    wire N__6374;
    wire N__6367;
    wire N__6364;
    wire N__6363;
    wire N__6360;
    wire N__6359;
    wire N__6356;
    wire N__6353;
    wire N__6350;
    wire N__6349;
    wire N__6346;
    wire N__6341;
    wire N__6338;
    wire N__6331;
    wire N__6330;
    wire N__6327;
    wire N__6324;
    wire N__6321;
    wire N__6320;
    wire N__6317;
    wire N__6316;
    wire N__6313;
    wire N__6310;
    wire N__6307;
    wire N__6304;
    wire N__6301;
    wire N__6298;
    wire N__6295;
    wire N__6292;
    wire N__6289;
    wire N__6286;
    wire N__6281;
    wire N__6274;
    wire N__6273;
    wire N__6272;
    wire N__6269;
    wire N__6266;
    wire N__6265;
    wire N__6262;
    wire N__6259;
    wire N__6256;
    wire N__6253;
    wire N__6250;
    wire N__6247;
    wire N__6244;
    wire N__6239;
    wire N__6236;
    wire N__6229;
    wire N__6228;
    wire N__6225;
    wire N__6222;
    wire N__6219;
    wire N__6216;
    wire N__6215;
    wire N__6210;
    wire N__6207;
    wire N__6204;
    wire N__6199;
    wire N__6196;
    wire N__6195;
    wire N__6194;
    wire N__6191;
    wire N__6188;
    wire N__6185;
    wire N__6178;
    wire N__6177;
    wire N__6174;
    wire N__6171;
    wire N__6170;
    wire N__6165;
    wire N__6162;
    wire N__6159;
    wire N__6156;
    wire N__6153;
    wire N__6150;
    wire N__6145;
    wire N__6142;
    wire N__6141;
    wire N__6138;
    wire N__6135;
    wire N__6132;
    wire N__6129;
    wire N__6128;
    wire N__6123;
    wire N__6120;
    wire N__6115;
    wire N__6114;
    wire N__6111;
    wire N__6108;
    wire N__6105;
    wire N__6102;
    wire N__6101;
    wire N__6100;
    wire N__6097;
    wire N__6094;
    wire N__6091;
    wire N__6088;
    wire N__6079;
    wire N__6078;
    wire N__6075;
    wire N__6074;
    wire N__6071;
    wire N__6070;
    wire N__6067;
    wire N__6064;
    wire N__6061;
    wire N__6058;
    wire N__6053;
    wire N__6050;
    wire N__6047;
    wire N__6044;
    wire N__6039;
    wire N__6036;
    wire N__6031;
    wire N__6030;
    wire N__6029;
    wire N__6028;
    wire N__6025;
    wire N__6022;
    wire N__6019;
    wire N__6016;
    wire N__6013;
    wire N__6010;
    wire N__6007;
    wire N__6004;
    wire N__6001;
    wire N__5994;
    wire N__5991;
    wire N__5988;
    wire N__5983;
    wire N__5980;
    wire N__5979;
    wire N__5976;
    wire N__5973;
    wire N__5970;
    wire N__5967;
    wire N__5966;
    wire N__5961;
    wire N__5958;
    wire N__5953;
    wire N__5950;
    wire N__5949;
    wire N__5948;
    wire N__5947;
    wire N__5946;
    wire N__5943;
    wire N__5940;
    wire N__5933;
    wire N__5930;
    wire N__5925;
    wire N__5920;
    wire N__5917;
    wire N__5914;
    wire N__5913;
    wire N__5910;
    wire N__5907;
    wire N__5906;
    wire N__5905;
    wire N__5902;
    wire N__5899;
    wire N__5896;
    wire N__5893;
    wire N__5884;
    wire N__5883;
    wire N__5880;
    wire N__5879;
    wire N__5878;
    wire N__5877;
    wire N__5874;
    wire N__5871;
    wire N__5864;
    wire N__5861;
    wire N__5856;
    wire N__5853;
    wire N__5848;
    wire N__5845;
    wire N__5842;
    wire N__5841;
    wire N__5838;
    wire N__5837;
    wire N__5834;
    wire N__5833;
    wire N__5830;
    wire N__5827;
    wire N__5824;
    wire N__5821;
    wire N__5816;
    wire N__5813;
    wire N__5810;
    wire N__5807;
    wire N__5802;
    wire N__5797;
    wire N__5794;
    wire N__5793;
    wire N__5792;
    wire N__5789;
    wire N__5786;
    wire N__5783;
    wire N__5780;
    wire N__5777;
    wire N__5774;
    wire N__5767;
    wire N__5764;
    wire N__5763;
    wire N__5760;
    wire N__5757;
    wire N__5754;
    wire N__5751;
    wire N__5750;
    wire N__5749;
    wire N__5748;
    wire N__5745;
    wire N__5742;
    wire N__5739;
    wire N__5736;
    wire N__5733;
    wire N__5730;
    wire N__5725;
    wire N__5720;
    wire N__5713;
    wire N__5710;
    wire N__5709;
    wire N__5706;
    wire N__5703;
    wire N__5702;
    wire N__5701;
    wire N__5700;
    wire N__5697;
    wire N__5694;
    wire N__5687;
    wire N__5680;
    wire N__5677;
    wire N__5674;
    wire N__5671;
    wire N__5668;
    wire N__5665;
    wire N__5662;
    wire N__5659;
    wire N__5658;
    wire N__5657;
    wire N__5656;
    wire N__5655;
    wire N__5654;
    wire N__5653;
    wire N__5652;
    wire N__5651;
    wire N__5650;
    wire N__5649;
    wire N__5648;
    wire N__5647;
    wire N__5646;
    wire N__5645;
    wire N__5644;
    wire N__5643;
    wire N__5642;
    wire N__5641;
    wire N__5640;
    wire N__5639;
    wire N__5638;
    wire N__5637;
    wire N__5636;
    wire N__5635;
    wire N__5634;
    wire N__5633;
    wire N__5632;
    wire N__5631;
    wire N__5630;
    wire N__5629;
    wire N__5628;
    wire N__5627;
    wire N__5626;
    wire N__5625;
    wire N__5624;
    wire N__5623;
    wire N__5548;
    wire N__5545;
    wire N__5542;
    wire N__5539;
    wire N__5536;
    wire N__5533;
    wire N__5530;
    wire N__5527;
    wire N__5524;
    wire N__5521;
    wire N__5520;
    wire N__5517;
    wire N__5516;
    wire N__5513;
    wire N__5510;
    wire N__5507;
    wire N__5502;
    wire N__5499;
    wire N__5494;
    wire N__5491;
    wire N__5488;
    wire N__5485;
    wire N__5484;
    wire N__5481;
    wire N__5478;
    wire N__5475;
    wire N__5472;
    wire N__5467;
    wire N__5464;
    wire N__5461;
    wire N__5458;
    wire N__5455;
    wire N__5452;
    wire N__5451;
    wire N__5448;
    wire N__5445;
    wire N__5442;
    wire N__5439;
    wire N__5436;
    wire N__5433;
    wire N__5430;
    wire N__5427;
    wire N__5422;
    wire N__5421;
    wire N__5420;
    wire N__5419;
    wire N__5418;
    wire N__5417;
    wire N__5416;
    wire N__5415;
    wire N__5414;
    wire N__5413;
    wire N__5410;
    wire N__5407;
    wire N__5402;
    wire N__5395;
    wire N__5388;
    wire N__5377;
    wire N__5376;
    wire N__5373;
    wire N__5370;
    wire N__5367;
    wire N__5362;
    wire N__5359;
    wire N__5358;
    wire N__5357;
    wire N__5356;
    wire N__5353;
    wire N__5350;
    wire N__5349;
    wire N__5346;
    wire N__5343;
    wire N__5342;
    wire N__5341;
    wire N__5340;
    wire N__5339;
    wire N__5336;
    wire N__5331;
    wire N__5328;
    wire N__5325;
    wire N__5322;
    wire N__5315;
    wire N__5302;
    wire N__5301;
    wire N__5300;
    wire N__5299;
    wire N__5298;
    wire N__5297;
    wire N__5294;
    wire N__5289;
    wire N__5284;
    wire N__5283;
    wire N__5280;
    wire N__5277;
    wire N__5272;
    wire N__5269;
    wire N__5266;
    wire N__5261;
    wire N__5258;
    wire N__5255;
    wire N__5250;
    wire N__5245;
    wire N__5244;
    wire N__5243;
    wire N__5242;
    wire N__5241;
    wire N__5238;
    wire N__5237;
    wire N__5234;
    wire N__5231;
    wire N__5226;
    wire N__5221;
    wire N__5214;
    wire N__5209;
    wire N__5206;
    wire N__5203;
    wire N__5200;
    wire N__5197;
    wire N__5194;
    wire N__5193;
    wire N__5192;
    wire N__5189;
    wire N__5186;
    wire N__5183;
    wire N__5182;
    wire N__5181;
    wire N__5178;
    wire N__5175;
    wire N__5172;
    wire N__5171;
    wire N__5168;
    wire N__5165;
    wire N__5160;
    wire N__5157;
    wire N__5154;
    wire N__5149;
    wire N__5146;
    wire N__5143;
    wire N__5134;
    wire N__5131;
    wire N__5128;
    wire N__5125;
    wire N__5124;
    wire N__5121;
    wire N__5118;
    wire N__5113;
    wire N__5110;
    wire N__5107;
    wire N__5104;
    wire N__5101;
    wire N__5100;
    wire N__5099;
    wire N__5096;
    wire N__5093;
    wire N__5092;
    wire N__5089;
    wire N__5086;
    wire N__5083;
    wire N__5082;
    wire N__5081;
    wire N__5080;
    wire N__5077;
    wire N__5074;
    wire N__5069;
    wire N__5064;
    wire N__5061;
    wire N__5058;
    wire N__5047;
    wire N__5044;
    wire N__5041;
    wire N__5038;
    wire N__5035;
    wire N__5032;
    wire N__5029;
    wire N__5028;
    wire N__5025;
    wire N__5022;
    wire N__5021;
    wire N__5016;
    wire N__5013;
    wire N__5012;
    wire N__5009;
    wire N__5006;
    wire N__5003;
    wire N__4996;
    wire N__4993;
    wire N__4990;
    wire N__4989;
    wire N__4988;
    wire N__4983;
    wire N__4982;
    wire N__4981;
    wire N__4980;
    wire N__4979;
    wire N__4978;
    wire N__4977;
    wire N__4974;
    wire N__4971;
    wire N__4968;
    wire N__4965;
    wire N__4962;
    wire N__4959;
    wire N__4954;
    wire N__4951;
    wire N__4936;
    wire N__4933;
    wire N__4932;
    wire N__4931;
    wire N__4930;
    wire N__4929;
    wire N__4928;
    wire N__4925;
    wire N__4922;
    wire N__4917;
    wire N__4914;
    wire N__4911;
    wire N__4910;
    wire N__4909;
    wire N__4908;
    wire N__4907;
    wire N__4906;
    wire N__4901;
    wire N__4898;
    wire N__4893;
    wire N__4888;
    wire N__4881;
    wire N__4870;
    wire N__4869;
    wire N__4866;
    wire N__4865;
    wire N__4864;
    wire N__4863;
    wire N__4860;
    wire N__4857;
    wire N__4850;
    wire N__4843;
    wire N__4842;
    wire N__4841;
    wire N__4840;
    wire N__4839;
    wire N__4836;
    wire N__4833;
    wire N__4830;
    wire N__4827;
    wire N__4824;
    wire N__4813;
    wire N__4810;
    wire N__4807;
    wire N__4806;
    wire N__4805;
    wire N__4800;
    wire N__4797;
    wire N__4792;
    wire N__4789;
    wire N__4786;
    wire N__4783;
    wire N__4782;
    wire N__4779;
    wire N__4776;
    wire N__4771;
    wire N__4768;
    wire N__4767;
    wire N__4764;
    wire N__4761;
    wire N__4760;
    wire N__4759;
    wire N__4758;
    wire N__4757;
    wire N__4754;
    wire N__4751;
    wire N__4746;
    wire N__4743;
    wire N__4740;
    wire N__4739;
    wire N__4738;
    wire N__4737;
    wire N__4736;
    wire N__4733;
    wire N__4730;
    wire N__4727;
    wire N__4714;
    wire N__4705;
    wire N__4704;
    wire N__4703;
    wire N__4702;
    wire N__4701;
    wire N__4700;
    wire N__4697;
    wire N__4692;
    wire N__4689;
    wire N__4686;
    wire N__4685;
    wire N__4684;
    wire N__4681;
    wire N__4678;
    wire N__4677;
    wire N__4674;
    wire N__4671;
    wire N__4668;
    wire N__4663;
    wire N__4658;
    wire N__4655;
    wire N__4642;
    wire N__4641;
    wire N__4638;
    wire N__4635;
    wire N__4630;
    wire N__4627;
    wire N__4624;
    wire N__4621;
    wire N__4618;
    wire N__4615;
    wire N__4612;
    wire N__4609;
    wire N__4606;
    wire N__4603;
    wire N__4600;
    wire N__4597;
    wire N__4594;
    wire N__4591;
    wire N__4588;
    wire N__4585;
    wire N__4582;
    wire N__4581;
    wire N__4578;
    wire N__4575;
    wire N__4572;
    wire N__4569;
    wire N__4564;
    wire N__4561;
    wire N__4558;
    wire N__4555;
    wire N__4554;
    wire N__4551;
    wire N__4548;
    wire N__4545;
    wire N__4540;
    wire N__4537;
    wire N__4534;
    wire N__4531;
    wire N__4528;
    wire N__4525;
    wire N__4524;
    wire N__4521;
    wire N__4518;
    wire N__4515;
    wire N__4510;
    wire N__4507;
    wire N__4504;
    wire N__4501;
    wire N__4500;
    wire N__4499;
    wire N__4496;
    wire N__4493;
    wire N__4490;
    wire N__4487;
    wire N__4480;
    wire N__4479;
    wire N__4478;
    wire N__4475;
    wire N__4472;
    wire N__4469;
    wire N__4468;
    wire N__4467;
    wire N__4466;
    wire N__4463;
    wire N__4460;
    wire N__4457;
    wire N__4454;
    wire N__4451;
    wire N__4448;
    wire N__4443;
    wire N__4438;
    wire N__4435;
    wire N__4430;
    wire N__4423;
    wire N__4420;
    wire N__4419;
    wire N__4418;
    wire N__4417;
    wire N__4416;
    wire N__4415;
    wire N__4412;
    wire N__4409;
    wire N__4406;
    wire N__4401;
    wire N__4400;
    wire N__4399;
    wire N__4398;
    wire N__4397;
    wire N__4396;
    wire N__4393;
    wire N__4390;
    wire N__4385;
    wire N__4382;
    wire N__4371;
    wire N__4368;
    wire N__4357;
    wire N__4354;
    wire N__4351;
    wire N__4348;
    wire N__4345;
    wire N__4342;
    wire N__4341;
    wire N__4338;
    wire N__4335;
    wire N__4330;
    wire N__4327;
    wire N__4326;
    wire N__4321;
    wire N__4320;
    wire N__4317;
    wire N__4314;
    wire N__4309;
    wire N__4306;
    wire N__4303;
    wire N__4300;
    wire N__4297;
    wire N__4296;
    wire N__4293;
    wire N__4290;
    wire N__4285;
    wire N__4282;
    wire N__4279;
    wire N__4276;
    wire N__4273;
    wire N__4270;
    wire N__4267;
    wire N__4264;
    wire N__4261;
    wire N__4258;
    wire N__4255;
    wire N__4252;
    wire N__4249;
    wire N__4246;
    wire N__4243;
    wire N__4240;
    wire N__4239;
    wire N__4236;
    wire N__4233;
    wire N__4228;
    wire N__4225;
    wire N__4224;
    wire N__4223;
    wire N__4220;
    wire N__4215;
    wire N__4210;
    wire N__4207;
    wire N__4204;
    wire N__4201;
    wire N__4200;
    wire N__4195;
    wire N__4194;
    wire N__4191;
    wire N__4188;
    wire N__4183;
    wire N__4180;
    wire N__4177;
    wire N__4174;
    wire N__4171;
    wire N__4168;
    wire N__4165;
    wire N__4162;
    wire N__4159;
    wire N__4156;
    wire N__4153;
    wire N__4150;
    wire N__4147;
    wire N__4144;
    wire N__4143;
    wire N__4142;
    wire N__4139;
    wire N__4138;
    wire N__4137;
    wire N__4136;
    wire N__4135;
    wire N__4132;
    wire N__4129;
    wire N__4128;
    wire N__4127;
    wire N__4124;
    wire N__4121;
    wire N__4118;
    wire N__4117;
    wire N__4116;
    wire N__4113;
    wire N__4110;
    wire N__4107;
    wire N__4104;
    wire N__4103;
    wire N__4102;
    wire N__4101;
    wire N__4098;
    wire N__4095;
    wire N__4092;
    wire N__4087;
    wire N__4080;
    wire N__4073;
    wire N__4070;
    wire N__4067;
    wire N__4062;
    wire N__4045;
    wire N__4044;
    wire N__4043;
    wire N__4042;
    wire N__4039;
    wire N__4034;
    wire N__4031;
    wire N__4028;
    wire N__4025;
    wire N__4024;
    wire N__4023;
    wire N__4022;
    wire N__4021;
    wire N__4020;
    wire N__4019;
    wire N__4014;
    wire N__4011;
    wire N__4006;
    wire N__4003;
    wire N__3996;
    wire N__3985;
    wire N__3982;
    wire N__3979;
    wire N__3978;
    wire N__3975;
    wire N__3972;
    wire N__3969;
    wire N__3966;
    wire N__3961;
    wire N__3958;
    wire N__3955;
    wire N__3952;
    wire N__3949;
    wire N__3946;
    wire N__3943;
    wire N__3940;
    wire N__3937;
    wire N__3934;
    wire N__3931;
    wire N__3928;
    wire N__3925;
    wire N__3924;
    wire N__3923;
    wire N__3920;
    wire N__3915;
    wire N__3910;
    wire N__3907;
    wire N__3904;
    wire N__3901;
    wire N__3898;
    wire N__3895;
    wire N__3892;
    wire N__3891;
    wire N__3888;
    wire N__3885;
    wire N__3884;
    wire N__3883;
    wire N__3880;
    wire N__3877;
    wire N__3874;
    wire N__3871;
    wire N__3868;
    wire N__3863;
    wire N__3856;
    wire N__3855;
    wire N__3850;
    wire N__3849;
    wire N__3848;
    wire N__3847;
    wire N__3844;
    wire N__3841;
    wire N__3838;
    wire N__3835;
    wire N__3826;
    wire N__3823;
    wire N__3820;
    wire N__3817;
    wire N__3814;
    wire N__3811;
    wire N__3810;
    wire N__3807;
    wire N__3804;
    wire N__3803;
    wire N__3798;
    wire N__3797;
    wire N__3794;
    wire N__3791;
    wire N__3788;
    wire N__3785;
    wire N__3778;
    wire N__3777;
    wire N__3776;
    wire N__3771;
    wire N__3768;
    wire N__3765;
    wire N__3760;
    wire N__3757;
    wire N__3754;
    wire N__3751;
    wire N__3748;
    wire N__3745;
    wire N__3742;
    wire N__3739;
    wire N__3736;
    wire N__3733;
    wire N__3732;
    wire N__3731;
    wire N__3728;
    wire N__3725;
    wire N__3722;
    wire N__3719;
    wire N__3716;
    wire N__3709;
    wire N__3708;
    wire N__3703;
    wire N__3700;
    wire N__3697;
    wire N__3694;
    wire N__3691;
    wire N__3688;
    wire N__3685;
    wire N__3682;
    wire N__3679;
    wire N__3676;
    wire N__3673;
    wire N__3670;
    wire N__3667;
    wire N__3664;
    wire N__3661;
    wire N__3658;
    wire N__3655;
    wire N__3652;
    wire N__3649;
    wire N__3648;
    wire N__3645;
    wire N__3642;
    wire N__3639;
    wire N__3636;
    wire N__3631;
    wire N__3628;
    wire N__3627;
    wire N__3624;
    wire N__3621;
    wire N__3616;
    wire N__3613;
    wire N__3610;
    wire N__3607;
    wire N__3604;
    wire N__3601;
    wire N__3598;
    wire N__3595;
    wire N__3592;
    wire N__3589;
    wire N__3588;
    wire N__3585;
    wire N__3584;
    wire N__3581;
    wire N__3578;
    wire N__3573;
    wire N__3570;
    wire N__3565;
    wire N__3562;
    wire N__3559;
    wire N__3558;
    wire N__3557;
    wire N__3554;
    wire N__3553;
    wire N__3552;
    wire N__3551;
    wire N__3548;
    wire N__3545;
    wire N__3544;
    wire N__3541;
    wire N__3534;
    wire N__3531;
    wire N__3528;
    wire N__3525;
    wire N__3522;
    wire N__3517;
    wire N__3512;
    wire N__3507;
    wire N__3502;
    wire N__3499;
    wire N__3496;
    wire N__3493;
    wire N__3490;
    wire N__3487;
    wire N__3484;
    wire N__3481;
    wire N__3478;
    wire N__3475;
    wire N__3472;
    wire N__3469;
    wire N__3466;
    wire N__3463;
    wire N__3460;
    wire N__3457;
    wire N__3454;
    wire N__3451;
    wire N__3448;
    wire N__3445;
    wire N__3444;
    wire N__3439;
    wire N__3436;
    wire N__3433;
    wire N__3430;
    wire N__3427;
    wire N__3424;
    wire N__3421;
    wire N__3418;
    wire N__3415;
    wire N__3412;
    wire N__3409;
    wire N__3406;
    wire N__3403;
    wire N__3400;
    wire N__3397;
    wire N__3394;
    wire N__3391;
    wire N__3388;
    wire N__3385;
    wire N__3382;
    wire N__3379;
    wire N__3376;
    wire N__3373;
    wire N__3370;
    wire N__3367;
    wire N__3364;
    wire N__3361;
    wire N__3358;
    wire N__3355;
    wire N__3352;
    wire N__3349;
    wire N__3346;
    wire N__3343;
    wire N__3340;
    wire N__3337;
    wire N__3334;
    wire N__3331;
    wire N__3328;
    wire N__3325;
    wire N__3322;
    wire N__3319;
    wire N__3318;
    wire N__3315;
    wire N__3312;
    wire N__3309;
    wire N__3306;
    wire N__3301;
    wire N__3298;
    wire N__3295;
    wire N__3292;
    wire N__3289;
    wire N__3288;
    wire N__3285;
    wire N__3282;
    wire N__3277;
    wire N__3274;
    wire N__3271;
    wire N__3268;
    wire N__3265;
    wire N__3262;
    wire N__3259;
    wire N__3256;
    wire N__3253;
    wire N__3250;
    wire N__3247;
    wire N__3244;
    wire N__3241;
    wire N__3238;
    wire N__3235;
    wire N__3232;
    wire N__3229;
    wire N__3226;
    wire VCCG0;
    wire GNDG0;
    wire G_138;
    wire G_138_cascade_;
    wire \uut.buf_clk_1 ;
    wire \INVuut.b_reg.ff6.qC_net ;
    wire \INVuut.b_reg.ff7.qC_net ;
    wire \INVuut.acc.ff2.qC_net ;
    wire \uut.AR_BUF.out_1_1_iv_3_1Z0Z_0_cascade_ ;
    wire \uut.AR_BUF.out_1_1_ivZ0Z_0_cascade_ ;
    wire \uut.out_1_1_iv_2_cascade_ ;
    wire \INVuut.AR.ff2.qC_net ;
    wire \uut.ALU_main.N_47_cascade_ ;
    wire \uut.seq.un1_HLT_1_reti_cascade_ ;
    wire \uut.un1_HLT_0 ;
    wire \INVuut.seq.q_ret_1C_net ;
    wire \uut.ALU_main.N_46_cascade_ ;
    wire \uut.alu_out_m_5_cascade_ ;
    wire \uut.bus_5_cascade_ ;
    wire \uut.alu_out_m_7_cascade_ ;
    wire \INVuut.b_reg.ff8.qC_net ;
    wire \uut.acc_out_m_7_cascade_ ;
    wire \uut.bus_7_cascade_ ;
    wire \uut.N_1_0 ;
    wire LED5_c;
    wire \INVuut.out_reg.ff5.qC_net ;
    wire \uut.out_1_2_iv_3_cascade_ ;
    wire LED1_c;
    wire \INVuut.out_reg.ff1.qC_net ;
    wire \INVuut.acc.ff3.qC_net ;
    wire \uut.program_counter_m_2_cascade_ ;
    wire \uut.AR_BUF.N_8 ;
    wire \uut.program_counter_m_2 ;
    wire \uut.AR_BUF.g0_0_0Z0Z_1 ;
    wire \uut.out_1_0_ivdup_2_cascade_ ;
    wire \uut.ALU_main.N_43 ;
    wire \uut.ir_out_m_d_1 ;
    wire \uut.bus_6_cascade_ ;
    wire \uut.q_RNIDGA71_cascade_ ;
    wire \INVuut.b_reg.ff5.qC_net ;
    wire \uut.ALU_main.N_45_cascade_ ;
    wire \uut.alu_out_m_4_cascade_ ;
    wire \uut.data_1_2_ivdup_cascade_ ;
    wire \uut.N_4_0 ;
    wire \uut.data_1_2_iv_0 ;
    wire \uut.b_reg_out_4 ;
    wire \INVuut.IR.ff5.q_0_neC_net ;
    wire \uut.AR_BUF.out_1_0_iv_2Z0Z_0 ;
    wire \uut.ir_out_m_d_2_cascade_ ;
    wire \INVuut.seq.q_retC_net ;
    wire \uut.ALU_main.N_48 ;
    wire \uut.AR_BUF.out_1_0_iv_2_1Z0Z_1 ;
    wire \INVuut.IR.ff1.q_neC_net ;
    wire \uut.AR_BUF.g0_0_a5_0Z0Z_2_cascade_ ;
    wire \uut.AR_BUF.N_9 ;
    wire \uut.AR_BUF.g0_1_a10_3Z0Z_2 ;
    wire \uut.AR_BUF.g0_0_o5_0Z0Z_0 ;
    wire \uut.AR_BUF.g0_1_a10_3_cascade_ ;
    wire \uut.AR_BUF.N_7 ;
    wire \uut.AR_BUF.N_13_cascade_ ;
    wire \uut.AR_BUF.g0_1_0Z0Z_5_cascade_ ;
    wire \uut.AR_BUF.g0_1_0Z0Z_1 ;
    wire \uut.AR_out_1 ;
    wire \uut.AR_BUF.g0_1_0_4_0 ;
    wire \uut.ir_out_1 ;
    wire \uut.AR_BUF.N_10 ;
    wire \uut.AR_BUF.g0_1_0_0_0 ;
    wire \uut.ir_out_m_d_0 ;
    wire \uut.pc.N_4_i_1_cascade_ ;
    wire \uut.alu_out_m_2 ;
    wire \INVuut.b_reg.ff3.qC_net ;
    wire \uut.ALU_main.N_43_0_cascade_ ;
    wire \uut.T_1_fast_RNIVM0N3_0_cascade_ ;
    wire \uut.pc.N_11 ;
    wire \uut.seq.counter.T_2_rep1_RNI8TEZ0Z81_cascade_ ;
    wire \uut.seq.counter.un2_MAR_LD_cascade_ ;
    wire \uut.D_1_0_cascade_ ;
    wire \uut.seq.q_ret_RNI52E81Z0Z_0 ;
    wire \uut.T_2_rep1_RNI6BLF1_cascade_ ;
    wire \uut.un17_IR_OE_0 ;
    wire \uut.IR.ir_out_m_c_d_1_3_cascade_ ;
    wire \uut.ir_out_m_c_d_3_cascade_ ;
    wire \INVuut.IR.ff4.q_neC_net ;
    wire \uut.seq.counter.T_2_rep1_RNIGC8CZ0Z1 ;
    wire \uut.seq.un13_ACC_LD_xZ0Z1_cascade_ ;
    wire \uut.un1_HLT_1 ;
    wire \uut.N_5_0 ;
    wire \uut.bus_6 ;
    wire \INVuut.IR.ff7.q_ret_1_fastC_net ;
    wire \uut.bus_7 ;
    wire \uut.seq.D_2_0_x_cascade_ ;
    wire \uut.q_0_fast ;
    wire \uut.data_1_2_ivdup ;
    wire \INVuut.IR.ff5.q_0_rep1C_net ;
    wire \uut.seq.counter.un4_ACC_LD_cascade_ ;
    wire \uut.seq.counter.ACC_LD_0_0 ;
    wire \uut.N_2_0 ;
    wire \INVuut.seq.counter.T_1_fast_3C_net ;
    wire \uut.q_ret_1_fast_0 ;
    wire \uut.AR_BUF.g0_3Z0Z_3_cascade_ ;
    wire \INVuut.acc.ff1.qC_net ;
    wire \uut.AR_BUF.out_1_2_ivZ0Z_1 ;
    wire \uut.ir_out_7 ;
    wire \uut.ir_out_6 ;
    wire \uut.AR_BUF.g0_3_a10_1Z0Z_1 ;
    wire \uut.D_1_0 ;
    wire \uut.AR_BUF.g0_3_a10_0Z0Z_2_cascade_ ;
    wire \uut.AR_BUF.g0_3Z0Z_0 ;
    wire \uut.ir_out_m_c_d_0_cascade_ ;
    wire \uut.AR_BUF.out_1_2_ivZ0Z_2 ;
    wire \uut.AR_BUF.g0_1_a10_4Z0Z_1 ;
    wire \uut.AR_BUF.g0_3Z0Z_2_cascade_ ;
    wire \uut.AR_BUF.g0_3Z0Z_6_cascade_ ;
    wire \INVuut.AR.ff1.q_neC_net ;
    wire \uut.AR_out_0 ;
    wire \uut.T_1_RNIVVKI3_3 ;
    wire \uut.program_counter_m_0 ;
    wire \uut.pc.G_26_i_a4_5_sx_cascade_ ;
    wire \uut.pc.G_26_i_a4_5 ;
    wire \uut.ir_out_m_c_c_0 ;
    wire \uut.alu_out_m_0_0 ;
    wire \uut.alu_out_m_0 ;
    wire \INVuut.b_reg.ff4.qC_net ;
    wire \uut.pc.program_counter_4_a1_0_0_1_cascade_ ;
    wire \uut.pc.g2_0 ;
    wire \uut.pc.N_77_0 ;
    wire \uut.pc.g1_0_cascade_ ;
    wire \uut.pc.program_counter_0_1_1 ;
    wire \uut.S0_0_i ;
    wire bfn_9_12_0_;
    wire \uut.un1_A_cry_0_s ;
    wire \uut.ALU_main.un1_A_cry_0_c_THRU_CO ;
    wire \uut.ALU_main.un1_A_cry_0 ;
    wire \uut.ALU_main.un1_A_cry_1_c_RNI7KLZ0Z45 ;
    wire \uut.ALU_main.un1_A_cry_1 ;
    wire \uut.ALU_main.un1_A_axb_3_l_ofxZ0 ;
    wire \uut.ALU_main.un1_A_cry_2_cZ0 ;
    wire \uut.ALU_main.un1_A_axb_4_l_ofxZ0 ;
    wire \uut.ALU_main.un1_A_cry_3_c_RNIF4UZ0Z45 ;
    wire \uut.ALU_main.un1_A_cry_3 ;
    wire \uut.ALU_main.un1_A_cry_4_c_RNIJCZ0Z255 ;
    wire \uut.ALU_main.un1_A_cry_4 ;
    wire \uut.ALU_main.un1_A_cry_5_c_RNINKZ0Z655 ;
    wire \uut.ALU_main.un1_A_cry_5 ;
    wire \uut.ALU_main.un1_A_cry_6 ;
    wire bfn_9_13_0_;
    wire \uut.ALU_main.un1_A_cry_6_c_RNINIMNZ0Z4 ;
    wire \uut.ALU_main.un1_A_axb_1_l_ofxZ0 ;
    wire \uut.b_reg_out_6 ;
    wire \uut.ALU_main.un1_A_axb_6_l_ofxZ0 ;
    wire \uut.b_reg_out_5 ;
    wire \uut.ALU_main.un1_A_axb_5_l_ofxZ0 ;
    wire \uut.ALU_main.un1_A_axb_0_l_ofxZ0 ;
    wire \uut.b_reg_out_7 ;
    wire \uut.ALU_main.un1_A_axbZ0Z_7 ;
    wire \uut.b_reg_out_2 ;
    wire \uut.acc_out_2 ;
    wire \uut.un13_ACC_LD ;
    wire \uut.ALU_main.un1_A_axb_2_l_ofxZ0 ;
    wire \uut.seq.counter.T_2_rep1_RNIJDGJZ0_cascade_ ;
    wire \uut.seq.D_4 ;
    wire \uut.D_1_3_cascade_ ;
    wire \uut.un7_ACC_LD ;
    wire \uut.ir_out_4 ;
    wire \uut.seq.counter.T_1_fastZ0Z_3 ;
    wire \uut.seq.counter.T_4_cascade_ ;
    wire \uut.seq.counter.T_1_fast_RNI4JTR1_0Z0Z_0 ;
    wire \uut.T_2_rep1 ;
    wire \uut.seq.counter.T_2_rep1_RNIV9NUZ0 ;
    wire \uut.bus_5 ;
    wire \uut.q_0_fast_1 ;
    wire \uut.seq.counter.T_1_fastZ0Z_0 ;
    wire \INVuut.IR.ff6.q_0_fastC_net ;
    wire \uut.ir_out_fast_4 ;
    wire \uut.ir_out_5 ;
    wire \uut.q_ret_1_fast ;
    wire \uut.seq.counter.T_4 ;
    wire \uut.seq.un10_ACC_LD_xZ0Z1_cascade_ ;
    wire \uut.T_1_fast_RNI28LI1_0_cascade_ ;
    wire \uut.N_41 ;
    wire \uut.q_0_fast_0 ;
    wire \uut.seq.counter.T_fastZ0Z_2 ;
    wire \uut.seq.counter.T_fast_RNIH09PZ0Z_2_cascade_ ;
    wire \uut.ir_out_4_rep1 ;
    wire \uut.ir_out_0 ;
    wire \uut.acc_out_0 ;
    wire \uut.OUT_LD_cascade_ ;
    wire \uut.pc.G_26_i_a4_1 ;
    wire \uut.acc_out_1 ;
    wire \uut.ALU_main.ALU_Out_0Z0Z_1_cascade_ ;
    wire \uut.un1_A_cry_0_c_RNI3CH45 ;
    wire \INVuut.seq.counter.T_1_4C_net ;
    wire \uut.seq.counter.un2_MAR_LD ;
    wire \uut.pc.g1 ;
    wire \uut.pc.un1_inc_0_0_cascade_ ;
    wire \INVuut.seq.counter.T_1_1C_net ;
    wire \uut.un17_IR_OE ;
    wire \uut.PC_LD_0_0 ;
    wire \uut.PC_LD_0_0_cascade_ ;
    wire \uut.pc.un1_inc_0 ;
    wire \uut.pc.un1_inc_0_cascade_ ;
    wire \uut.pc.program_counter_4_1_2 ;
    wire \uut.m13 ;
    wire \INVuut.mar.ff2.q_neC_net ;
    wire \uut.program_counter_2 ;
    wire \uut.program_counter_1 ;
    wire \uut.program_counter_0 ;
    wire \uut.pc.program_counter_RNO_1Z0Z_2 ;
    wire \uut.N_44_0_cascade_ ;
    wire \uut.pc.g0_rn_1 ;
    wire \uut.pc.alu_out_m_0_3_cascade_ ;
    wire \uut.buf_clk_1_g ;
    wire \uut.ALU_main.N_44_1 ;
    wire \uut.T_1_fast_RNI28LI1_0 ;
    wire \uut.b_reg_out_3 ;
    wire \uut.un1_A_cry_2_c_RNIBSP45 ;
    wire \uut.un1_ALU_en_0 ;
    wire \uut.ALU_main.N_44_cascade_ ;
    wire \uut.T_1_fast_RNIVM0N3_0 ;
    wire \uut.acc_out_m_6 ;
    wire \uut.alu_out_m_6 ;
    wire \uut.mem.N_29_mux ;
    wire \uut.acc_out_6 ;
    wire \uut.acc_out_m_7 ;
    wire \uut.alu_out_m_7 ;
    wire \uut.acc_out_7 ;
    wire \uut.alu_out_m_5 ;
    wire \uut.acc_out_m_5 ;
    wire \uut.mem.m20 ;
    wire \uut.acc_out_5 ;
    wire \uut.q_RNIDGA71 ;
    wire \uut.mem.i2_mux ;
    wire \uut.alu_out_m_4 ;
    wire \uut.acc_out_4 ;
    wire \INVuut.acc.ff4.qC_net ;
    wire \uut.ACC_LD_0_i ;
    wire \uut.seq.D_2_1 ;
    wire \uut.ir_out_i_2_6 ;
    wire \uut.seq.D_2 ;
    wire \uut.ir_out_i_2_5 ;
    wire \uut.B_LD_0_1_tz_cascade_ ;
    wire \uut.mem.i2_mux_0 ;
    wire \uut.out_1_0_iv_2_1 ;
    wire LED3_c;
    wire \INVuut.out_reg.ff3.qC_net ;
    wire \uut.m10 ;
    wire \uut.m10_cascade_ ;
    wire \uut.b_reg_out_0 ;
    wire \uut.alu_out_m_1 ;
    wire \uut.N_11_i_m ;
    wire \uut.out_1_1_iv_3dup_1 ;
    wire \uut.b_reg_out_1 ;
    wire \INVuut.b_reg.ff1.qC_net ;
    wire \uut.B_LD_0_i ;
    wire \uut.inc ;
    wire \uut.ir_out_2 ;
    wire \INVuut.IR.ff3.qC_net ;
    wire \uut.N_14_0 ;
    wire \uut.alu_out_m_0_2 ;
    wire \uut.out_1_0_iv_3_cascade_ ;
    wire \uut.AR_out_2 ;
    wire \INVuut.AR.ff3.qC_net ;
    wire \uut.un11_MAR_LD ;
    wire \uut.MAR_LD_1 ;
    wire \uut.seq.counter.MAR_LD_0_0 ;
    wire \uut.MAR_LD_1_cascade_ ;
    wire \uut.N_16_0 ;
    wire \uut.alu_out_m_1_3 ;
    wire \uut.AR_BUF.g0Z0Z_5_cascade_ ;
    wire \INVuut.AR.ff4.q_neC_net ;
    wire \uut.AR_LD ;
    wire \uut.un14_MAR_LD ;
    wire \uut.un8_MAR_LD ;
    wire \uut.un1_IR_OE_4_1 ;
    wire \uut.pc.un1_inc_0_0 ;
    wire \uut.ir_out_m_d_3_cascade_ ;
    wire \uut.pc.g0_sn ;
    wire \uut.seq.counter.T_1Z0Z_4 ;
    wire \INVuut.seq.counter.T_1_0C_net ;
    wire \uut.AR_BUF.out_1_ivdupZ0Z_0_cascade_ ;
    wire \uut.g0_0 ;
    wire \uut.AR_out_3 ;
    wire \uut.g1_cascade_ ;
    wire \uut.T_2_rep1_RNI6BLF1 ;
    wire \uut.AR_BUF.g0_1_0 ;
    wire \uut.T_2 ;
    wire \uut.T_0 ;
    wire \uut.program_counter_3 ;
    wire \uut.D_6 ;
    wire \uut.program_counter_m_3 ;
    wire \uut.acc_out_3 ;
    wire \uut.ir_out_3 ;
    wire \uut.un5_MAR_LD ;
    wire \uut.AR_BUF.out_1_ivZ0Z_0_cascade_ ;
    wire \uut.out_1_iv_2 ;
    wire \uut.out_1_iv_2_1_cascade_ ;
    wire \uut.OUT_LD ;
    wire LED4_c;
    wire \uut.alu_out_m_3 ;
    wire \uut.m15_cascade_ ;
    wire \uut.out_1_iv_3 ;
    wire \uut.out_1_0_ivdup_2 ;
    wire \uut.out_1_0_iv_3 ;
    wire \uut.MAR_LD_0 ;
    wire \INVuut.out_reg.ff4.qC_net ;
    wire \uut.g1_0 ;
    wire \uut.ir_out_m_d_3 ;
    wire \uut.AR_BUF.g0Z0Z_5 ;
    wire \uut.AR_BUF.g0_0Z0Z_0 ;
    wire \uut.ir_out_m_c_d_3 ;
    wire \uut.mar_out_2 ;
    wire \uut.mar_out_3 ;
    wire \uut.mar_out_1 ;
    wire \uut.seq.counter.T_1_fast_RNI6J9SZ0Z_3 ;
    wire \uut.D_1_3 ;
    wire \uut.seq.counter.T_1_fastZ0Z_1 ;
    wire \uut.T_3 ;
    wire \uut.un1_ROM_OE_0_cascade_ ;
    wire \uut.B_LD_0_1_tz ;
    wire \uut.un1_ROM_OE_0 ;
    wire \uut.mem.N_7_i_m_sx_cascade_ ;
    wire \uut.B_LD_0_2_tz ;
    wire \uut.N_7_i_m ;
    wire \uut.AR_BUF.g0_3Z0Z_6 ;
    wire \uut.AR_BUF.g0_3Z0Z_3 ;
    wire \uut.m6 ;
    wire \uut.ROM_OE ;
    wire \uut.mar_out_0 ;
    wire \INVuut.mar.ff4.q_neC_net ;
    wire \uut.mar.MAR_LD_0_1 ;
    wire _gnd_net_;

    defparam LED1_obuf_iopad.PULLUP=1'b0;
    defparam LED1_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD LED1_obuf_iopad (
            .OE(N__9920),
            .DIN(N__9919),
            .DOUT(N__9918),
            .PACKAGEPIN(LED1));
    defparam LED1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED1_obuf_preio (
            .PADOEN(N__9920),
            .PADOUT(N__9919),
            .PADIN(N__9918),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3298),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam LED4_obuf_iopad.PULLUP=1'b0;
    defparam LED4_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD LED4_obuf_iopad (
            .OE(N__9911),
            .DIN(N__9910),
            .DOUT(N__9909),
            .PACKAGEPIN(LED4));
    defparam LED4_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED4_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED4_obuf_preio (
            .PADOEN(N__9911),
            .PADOUT(N__9910),
            .PADIN(N__9909),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__8161),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam LED2_obuf_iopad.PULLUP=1'b0;
    defparam LED2_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD LED2_obuf_iopad (
            .OE(N__9902),
            .DIN(N__9901),
            .DOUT(N__9900),
            .PACKAGEPIN(LED2));
    defparam LED2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED2_obuf_preio (
            .PADOEN(N__9902),
            .PADOUT(N__9901),
            .PADIN(N__9900),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(GNDG0),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam LED3_obuf_iopad.PULLUP=1'b0;
    defparam LED3_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD LED3_obuf_iopad (
            .OE(N__9893),
            .DIN(N__9892),
            .DOUT(N__9891),
            .PACKAGEPIN(LED3));
    defparam LED3_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED3_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED3_obuf_preio (
            .PADOEN(N__9893),
            .PADOUT(N__9892),
            .PADIN(N__9891),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__6838),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    defparam LED5_obuf_iopad.PULLUP=1'b0;
    defparam LED5_obuf_iopad.IO_STANDARD="SB_LVCMOS";
    IO_PAD LED5_obuf_iopad (
            .OE(N__9884),
            .DIN(N__9883),
            .DOUT(N__9882),
            .PACKAGEPIN(LED5));
    defparam LED5_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED5_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED5_obuf_preio (
            .PADOEN(N__9884),
            .PADOUT(N__9883),
            .PADIN(N__9882),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__3328),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    InMux I__2509 (
            .O(N__9865),
            .I(N__9862));
    LocalMux I__2508 (
            .O(N__9862),
            .I(\uut.g1_0 ));
    InMux I__2507 (
            .O(N__9859),
            .I(N__9856));
    LocalMux I__2506 (
            .O(N__9856),
            .I(N__9853));
    Span4Mux_v I__2505 (
            .O(N__9853),
            .I(N__9847));
    InMux I__2504 (
            .O(N__9852),
            .I(N__9844));
    InMux I__2503 (
            .O(N__9851),
            .I(N__9841));
    InMux I__2502 (
            .O(N__9850),
            .I(N__9837));
    Span4Mux_h I__2501 (
            .O(N__9847),
            .I(N__9829));
    LocalMux I__2500 (
            .O(N__9844),
            .I(N__9829));
    LocalMux I__2499 (
            .O(N__9841),
            .I(N__9829));
    InMux I__2498 (
            .O(N__9840),
            .I(N__9826));
    LocalMux I__2497 (
            .O(N__9837),
            .I(N__9823));
    InMux I__2496 (
            .O(N__9836),
            .I(N__9820));
    Sp12to4 I__2495 (
            .O(N__9829),
            .I(N__9815));
    LocalMux I__2494 (
            .O(N__9826),
            .I(N__9815));
    Odrv4 I__2493 (
            .O(N__9823),
            .I(\uut.ir_out_m_d_3 ));
    LocalMux I__2492 (
            .O(N__9820),
            .I(\uut.ir_out_m_d_3 ));
    Odrv12 I__2491 (
            .O(N__9815),
            .I(\uut.ir_out_m_d_3 ));
    InMux I__2490 (
            .O(N__9808),
            .I(N__9805));
    LocalMux I__2489 (
            .O(N__9805),
            .I(N__9799));
    InMux I__2488 (
            .O(N__9804),
            .I(N__9796));
    InMux I__2487 (
            .O(N__9803),
            .I(N__9793));
    InMux I__2486 (
            .O(N__9802),
            .I(N__9790));
    Span4Mux_h I__2485 (
            .O(N__9799),
            .I(N__9785));
    LocalMux I__2484 (
            .O(N__9796),
            .I(N__9785));
    LocalMux I__2483 (
            .O(N__9793),
            .I(N__9782));
    LocalMux I__2482 (
            .O(N__9790),
            .I(N__9779));
    Odrv4 I__2481 (
            .O(N__9785),
            .I(\uut.AR_BUF.g0Z0Z_5 ));
    Odrv12 I__2480 (
            .O(N__9782),
            .I(\uut.AR_BUF.g0Z0Z_5 ));
    Odrv12 I__2479 (
            .O(N__9779),
            .I(\uut.AR_BUF.g0Z0Z_5 ));
    CascadeMux I__2478 (
            .O(N__9772),
            .I(N__9768));
    CascadeMux I__2477 (
            .O(N__9771),
            .I(N__9764));
    InMux I__2476 (
            .O(N__9768),
            .I(N__9760));
    InMux I__2475 (
            .O(N__9767),
            .I(N__9757));
    InMux I__2474 (
            .O(N__9764),
            .I(N__9754));
    CascadeMux I__2473 (
            .O(N__9763),
            .I(N__9751));
    LocalMux I__2472 (
            .O(N__9760),
            .I(N__9748));
    LocalMux I__2471 (
            .O(N__9757),
            .I(N__9743));
    LocalMux I__2470 (
            .O(N__9754),
            .I(N__9743));
    InMux I__2469 (
            .O(N__9751),
            .I(N__9740));
    Span4Mux_s3_h I__2468 (
            .O(N__9748),
            .I(N__9736));
    Span4Mux_s3_h I__2467 (
            .O(N__9743),
            .I(N__9733));
    LocalMux I__2466 (
            .O(N__9740),
            .I(N__9730));
    InMux I__2465 (
            .O(N__9739),
            .I(N__9727));
    Odrv4 I__2464 (
            .O(N__9736),
            .I(\uut.AR_BUF.g0_0Z0Z_0 ));
    Odrv4 I__2463 (
            .O(N__9733),
            .I(\uut.AR_BUF.g0_0Z0Z_0 ));
    Odrv4 I__2462 (
            .O(N__9730),
            .I(\uut.AR_BUF.g0_0Z0Z_0 ));
    LocalMux I__2461 (
            .O(N__9727),
            .I(\uut.AR_BUF.g0_0Z0Z_0 ));
    InMux I__2460 (
            .O(N__9718),
            .I(N__9715));
    LocalMux I__2459 (
            .O(N__9715),
            .I(N__9708));
    InMux I__2458 (
            .O(N__9714),
            .I(N__9705));
    InMux I__2457 (
            .O(N__9713),
            .I(N__9702));
    InMux I__2456 (
            .O(N__9712),
            .I(N__9697));
    InMux I__2455 (
            .O(N__9711),
            .I(N__9697));
    Span4Mux_v I__2454 (
            .O(N__9708),
            .I(N__9692));
    LocalMux I__2453 (
            .O(N__9705),
            .I(N__9692));
    LocalMux I__2452 (
            .O(N__9702),
            .I(N__9687));
    LocalMux I__2451 (
            .O(N__9697),
            .I(N__9687));
    Span4Mux_s3_v I__2450 (
            .O(N__9692),
            .I(N__9684));
    Span12Mux_s4_h I__2449 (
            .O(N__9687),
            .I(N__9681));
    Odrv4 I__2448 (
            .O(N__9684),
            .I(\uut.ir_out_m_c_d_3 ));
    Odrv12 I__2447 (
            .O(N__9681),
            .I(\uut.ir_out_m_c_d_3 ));
    CascadeMux I__2446 (
            .O(N__9676),
            .I(N__9672));
    CascadeMux I__2445 (
            .O(N__9675),
            .I(N__9667));
    InMux I__2444 (
            .O(N__9672),
            .I(N__9656));
    InMux I__2443 (
            .O(N__9671),
            .I(N__9656));
    InMux I__2442 (
            .O(N__9670),
            .I(N__9656));
    InMux I__2441 (
            .O(N__9667),
            .I(N__9656));
    InMux I__2440 (
            .O(N__9666),
            .I(N__9645));
    InMux I__2439 (
            .O(N__9665),
            .I(N__9645));
    LocalMux I__2438 (
            .O(N__9656),
            .I(N__9642));
    InMux I__2437 (
            .O(N__9655),
            .I(N__9637));
    InMux I__2436 (
            .O(N__9654),
            .I(N__9637));
    InMux I__2435 (
            .O(N__9653),
            .I(N__9632));
    InMux I__2434 (
            .O(N__9652),
            .I(N__9632));
    InMux I__2433 (
            .O(N__9651),
            .I(N__9629));
    InMux I__2432 (
            .O(N__9650),
            .I(N__9626));
    LocalMux I__2431 (
            .O(N__9645),
            .I(\uut.mar_out_2 ));
    Odrv4 I__2430 (
            .O(N__9642),
            .I(\uut.mar_out_2 ));
    LocalMux I__2429 (
            .O(N__9637),
            .I(\uut.mar_out_2 ));
    LocalMux I__2428 (
            .O(N__9632),
            .I(\uut.mar_out_2 ));
    LocalMux I__2427 (
            .O(N__9629),
            .I(\uut.mar_out_2 ));
    LocalMux I__2426 (
            .O(N__9626),
            .I(\uut.mar_out_2 ));
    CascadeMux I__2425 (
            .O(N__9613),
            .I(N__9604));
    CascadeMux I__2424 (
            .O(N__9612),
            .I(N__9601));
    CascadeMux I__2423 (
            .O(N__9611),
            .I(N__9597));
    CascadeMux I__2422 (
            .O(N__9610),
            .I(N__9594));
    CascadeMux I__2421 (
            .O(N__9609),
            .I(N__9591));
    CascadeMux I__2420 (
            .O(N__9608),
            .I(N__9586));
    InMux I__2419 (
            .O(N__9607),
            .I(N__9577));
    InMux I__2418 (
            .O(N__9604),
            .I(N__9577));
    InMux I__2417 (
            .O(N__9601),
            .I(N__9577));
    InMux I__2416 (
            .O(N__9600),
            .I(N__9577));
    InMux I__2415 (
            .O(N__9597),
            .I(N__9572));
    InMux I__2414 (
            .O(N__9594),
            .I(N__9572));
    InMux I__2413 (
            .O(N__9591),
            .I(N__9566));
    InMux I__2412 (
            .O(N__9590),
            .I(N__9566));
    InMux I__2411 (
            .O(N__9589),
            .I(N__9561));
    InMux I__2410 (
            .O(N__9586),
            .I(N__9561));
    LocalMux I__2409 (
            .O(N__9577),
            .I(N__9556));
    LocalMux I__2408 (
            .O(N__9572),
            .I(N__9556));
    InMux I__2407 (
            .O(N__9571),
            .I(N__9553));
    LocalMux I__2406 (
            .O(N__9566),
            .I(\uut.mar_out_3 ));
    LocalMux I__2405 (
            .O(N__9561),
            .I(\uut.mar_out_3 ));
    Odrv4 I__2404 (
            .O(N__9556),
            .I(\uut.mar_out_3 ));
    LocalMux I__2403 (
            .O(N__9553),
            .I(\uut.mar_out_3 ));
    CascadeMux I__2402 (
            .O(N__9544),
            .I(N__9540));
    CascadeMux I__2401 (
            .O(N__9543),
            .I(N__9536));
    InMux I__2400 (
            .O(N__9540),
            .I(N__9530));
    InMux I__2399 (
            .O(N__9539),
            .I(N__9530));
    InMux I__2398 (
            .O(N__9536),
            .I(N__9527));
    InMux I__2397 (
            .O(N__9535),
            .I(N__9517));
    LocalMux I__2396 (
            .O(N__9530),
            .I(N__9512));
    LocalMux I__2395 (
            .O(N__9527),
            .I(N__9512));
    InMux I__2394 (
            .O(N__9526),
            .I(N__9509));
    InMux I__2393 (
            .O(N__9525),
            .I(N__9500));
    InMux I__2392 (
            .O(N__9524),
            .I(N__9500));
    InMux I__2391 (
            .O(N__9523),
            .I(N__9500));
    InMux I__2390 (
            .O(N__9522),
            .I(N__9500));
    InMux I__2389 (
            .O(N__9521),
            .I(N__9495));
    InMux I__2388 (
            .O(N__9520),
            .I(N__9495));
    LocalMux I__2387 (
            .O(N__9517),
            .I(N__9490));
    Span4Mux_s3_v I__2386 (
            .O(N__9512),
            .I(N__9490));
    LocalMux I__2385 (
            .O(N__9509),
            .I(\uut.mar_out_1 ));
    LocalMux I__2384 (
            .O(N__9500),
            .I(\uut.mar_out_1 ));
    LocalMux I__2383 (
            .O(N__9495),
            .I(\uut.mar_out_1 ));
    Odrv4 I__2382 (
            .O(N__9490),
            .I(\uut.mar_out_1 ));
    InMux I__2381 (
            .O(N__9481),
            .I(N__9478));
    LocalMux I__2380 (
            .O(N__9478),
            .I(N__9475));
    Span4Mux_s3_h I__2379 (
            .O(N__9475),
            .I(N__9472));
    Odrv4 I__2378 (
            .O(N__9472),
            .I(\uut.seq.counter.T_1_fast_RNI6J9SZ0Z_3 ));
    InMux I__2377 (
            .O(N__9469),
            .I(N__9465));
    InMux I__2376 (
            .O(N__9468),
            .I(N__9461));
    LocalMux I__2375 (
            .O(N__9465),
            .I(N__9455));
    InMux I__2374 (
            .O(N__9464),
            .I(N__9452));
    LocalMux I__2373 (
            .O(N__9461),
            .I(N__9449));
    InMux I__2372 (
            .O(N__9460),
            .I(N__9446));
    InMux I__2371 (
            .O(N__9459),
            .I(N__9441));
    InMux I__2370 (
            .O(N__9458),
            .I(N__9441));
    Span4Mux_s2_v I__2369 (
            .O(N__9455),
            .I(N__9436));
    LocalMux I__2368 (
            .O(N__9452),
            .I(N__9436));
    Odrv12 I__2367 (
            .O(N__9449),
            .I(\uut.D_1_3 ));
    LocalMux I__2366 (
            .O(N__9446),
            .I(\uut.D_1_3 ));
    LocalMux I__2365 (
            .O(N__9441),
            .I(\uut.D_1_3 ));
    Odrv4 I__2364 (
            .O(N__9436),
            .I(\uut.D_1_3 ));
    InMux I__2363 (
            .O(N__9427),
            .I(N__9424));
    LocalMux I__2362 (
            .O(N__9424),
            .I(N__9421));
    Span4Mux_s2_h I__2361 (
            .O(N__9421),
            .I(N__9416));
    InMux I__2360 (
            .O(N__9420),
            .I(N__9413));
    InMux I__2359 (
            .O(N__9419),
            .I(N__9410));
    Odrv4 I__2358 (
            .O(N__9416),
            .I(\uut.seq.counter.T_1_fastZ0Z_1 ));
    LocalMux I__2357 (
            .O(N__9413),
            .I(\uut.seq.counter.T_1_fastZ0Z_1 ));
    LocalMux I__2356 (
            .O(N__9410),
            .I(\uut.seq.counter.T_1_fastZ0Z_1 ));
    InMux I__2355 (
            .O(N__9403),
            .I(N__9397));
    InMux I__2354 (
            .O(N__9402),
            .I(N__9390));
    InMux I__2353 (
            .O(N__9401),
            .I(N__9387));
    InMux I__2352 (
            .O(N__9400),
            .I(N__9384));
    LocalMux I__2351 (
            .O(N__9397),
            .I(N__9381));
    InMux I__2350 (
            .O(N__9396),
            .I(N__9378));
    InMux I__2349 (
            .O(N__9395),
            .I(N__9373));
    InMux I__2348 (
            .O(N__9394),
            .I(N__9373));
    InMux I__2347 (
            .O(N__9393),
            .I(N__9370));
    LocalMux I__2346 (
            .O(N__9390),
            .I(N__9367));
    LocalMux I__2345 (
            .O(N__9387),
            .I(N__9364));
    LocalMux I__2344 (
            .O(N__9384),
            .I(N__9357));
    Span4Mux_h I__2343 (
            .O(N__9381),
            .I(N__9357));
    LocalMux I__2342 (
            .O(N__9378),
            .I(N__9353));
    LocalMux I__2341 (
            .O(N__9373),
            .I(N__9350));
    LocalMux I__2340 (
            .O(N__9370),
            .I(N__9345));
    Span4Mux_h I__2339 (
            .O(N__9367),
            .I(N__9345));
    Span4Mux_h I__2338 (
            .O(N__9364),
            .I(N__9342));
    InMux I__2337 (
            .O(N__9363),
            .I(N__9337));
    InMux I__2336 (
            .O(N__9362),
            .I(N__9337));
    Span4Mux_v I__2335 (
            .O(N__9357),
            .I(N__9334));
    InMux I__2334 (
            .O(N__9356),
            .I(N__9331));
    Span4Mux_h I__2333 (
            .O(N__9353),
            .I(N__9324));
    Span4Mux_h I__2332 (
            .O(N__9350),
            .I(N__9324));
    Span4Mux_v I__2331 (
            .O(N__9345),
            .I(N__9324));
    Odrv4 I__2330 (
            .O(N__9342),
            .I(\uut.T_3 ));
    LocalMux I__2329 (
            .O(N__9337),
            .I(\uut.T_3 ));
    Odrv4 I__2328 (
            .O(N__9334),
            .I(\uut.T_3 ));
    LocalMux I__2327 (
            .O(N__9331),
            .I(\uut.T_3 ));
    Odrv4 I__2326 (
            .O(N__9324),
            .I(\uut.T_3 ));
    CascadeMux I__2325 (
            .O(N__9313),
            .I(\uut.un1_ROM_OE_0_cascade_ ));
    InMux I__2324 (
            .O(N__9310),
            .I(N__9306));
    InMux I__2323 (
            .O(N__9309),
            .I(N__9303));
    LocalMux I__2322 (
            .O(N__9306),
            .I(\uut.B_LD_0_1_tz ));
    LocalMux I__2321 (
            .O(N__9303),
            .I(\uut.B_LD_0_1_tz ));
    InMux I__2320 (
            .O(N__9298),
            .I(N__9294));
    InMux I__2319 (
            .O(N__9297),
            .I(N__9291));
    LocalMux I__2318 (
            .O(N__9294),
            .I(\uut.un1_ROM_OE_0 ));
    LocalMux I__2317 (
            .O(N__9291),
            .I(\uut.un1_ROM_OE_0 ));
    CascadeMux I__2316 (
            .O(N__9286),
            .I(\uut.mem.N_7_i_m_sx_cascade_ ));
    InMux I__2315 (
            .O(N__9283),
            .I(N__9280));
    LocalMux I__2314 (
            .O(N__9280),
            .I(N__9275));
    InMux I__2313 (
            .O(N__9279),
            .I(N__9270));
    InMux I__2312 (
            .O(N__9278),
            .I(N__9270));
    Span4Mux_s0_h I__2311 (
            .O(N__9275),
            .I(N__9265));
    LocalMux I__2310 (
            .O(N__9270),
            .I(N__9265));
    Odrv4 I__2309 (
            .O(N__9265),
            .I(\uut.B_LD_0_2_tz ));
    InMux I__2308 (
            .O(N__9262),
            .I(N__9259));
    LocalMux I__2307 (
            .O(N__9259),
            .I(N__9255));
    InMux I__2306 (
            .O(N__9258),
            .I(N__9252));
    Span4Mux_v I__2305 (
            .O(N__9255),
            .I(N__9247));
    LocalMux I__2304 (
            .O(N__9252),
            .I(N__9247));
    Span4Mux_h I__2303 (
            .O(N__9247),
            .I(N__9244));
    Odrv4 I__2302 (
            .O(N__9244),
            .I(\uut.N_7_i_m ));
    InMux I__2301 (
            .O(N__9241),
            .I(N__9236));
    InMux I__2300 (
            .O(N__9240),
            .I(N__9233));
    InMux I__2299 (
            .O(N__9239),
            .I(N__9230));
    LocalMux I__2298 (
            .O(N__9236),
            .I(N__9227));
    LocalMux I__2297 (
            .O(N__9233),
            .I(N__9224));
    LocalMux I__2296 (
            .O(N__9230),
            .I(N__9221));
    Span4Mux_s2_h I__2295 (
            .O(N__9227),
            .I(N__9217));
    Span4Mux_s3_h I__2294 (
            .O(N__9224),
            .I(N__9212));
    Span4Mux_h I__2293 (
            .O(N__9221),
            .I(N__9212));
    InMux I__2292 (
            .O(N__9220),
            .I(N__9209));
    Span4Mux_v I__2291 (
            .O(N__9217),
            .I(N__9206));
    Span4Mux_v I__2290 (
            .O(N__9212),
            .I(N__9201));
    LocalMux I__2289 (
            .O(N__9209),
            .I(N__9201));
    Odrv4 I__2288 (
            .O(N__9206),
            .I(\uut.AR_BUF.g0_3Z0Z_6 ));
    Odrv4 I__2287 (
            .O(N__9201),
            .I(\uut.AR_BUF.g0_3Z0Z_6 ));
    InMux I__2286 (
            .O(N__9196),
            .I(N__9191));
    CascadeMux I__2285 (
            .O(N__9195),
            .I(N__9188));
    CascadeMux I__2284 (
            .O(N__9194),
            .I(N__9185));
    LocalMux I__2283 (
            .O(N__9191),
            .I(N__9182));
    InMux I__2282 (
            .O(N__9188),
            .I(N__9179));
    InMux I__2281 (
            .O(N__9185),
            .I(N__9176));
    Span4Mux_v I__2280 (
            .O(N__9182),
            .I(N__9172));
    LocalMux I__2279 (
            .O(N__9179),
            .I(N__9169));
    LocalMux I__2278 (
            .O(N__9176),
            .I(N__9166));
    InMux I__2277 (
            .O(N__9175),
            .I(N__9163));
    Span4Mux_h I__2276 (
            .O(N__9172),
            .I(N__9158));
    Span4Mux_v I__2275 (
            .O(N__9169),
            .I(N__9158));
    Span4Mux_v I__2274 (
            .O(N__9166),
            .I(N__9155));
    LocalMux I__2273 (
            .O(N__9163),
            .I(N__9152));
    Span4Mux_v I__2272 (
            .O(N__9158),
            .I(N__9147));
    Span4Mux_v I__2271 (
            .O(N__9155),
            .I(N__9147));
    Span4Mux_v I__2270 (
            .O(N__9152),
            .I(N__9144));
    Odrv4 I__2269 (
            .O(N__9147),
            .I(\uut.AR_BUF.g0_3Z0Z_3 ));
    Odrv4 I__2268 (
            .O(N__9144),
            .I(\uut.AR_BUF.g0_3Z0Z_3 ));
    InMux I__2267 (
            .O(N__9139),
            .I(N__9134));
    InMux I__2266 (
            .O(N__9138),
            .I(N__9130));
    InMux I__2265 (
            .O(N__9137),
            .I(N__9127));
    LocalMux I__2264 (
            .O(N__9134),
            .I(N__9124));
    CascadeMux I__2263 (
            .O(N__9133),
            .I(N__9120));
    LocalMux I__2262 (
            .O(N__9130),
            .I(N__9117));
    LocalMux I__2261 (
            .O(N__9127),
            .I(N__9114));
    Span4Mux_h I__2260 (
            .O(N__9124),
            .I(N__9111));
    InMux I__2259 (
            .O(N__9123),
            .I(N__9107));
    InMux I__2258 (
            .O(N__9120),
            .I(N__9104));
    Span4Mux_h I__2257 (
            .O(N__9117),
            .I(N__9101));
    Span12Mux_s2_v I__2256 (
            .O(N__9114),
            .I(N__9098));
    Span4Mux_v I__2255 (
            .O(N__9111),
            .I(N__9095));
    InMux I__2254 (
            .O(N__9110),
            .I(N__9092));
    LocalMux I__2253 (
            .O(N__9107),
            .I(\uut.m6 ));
    LocalMux I__2252 (
            .O(N__9104),
            .I(\uut.m6 ));
    Odrv4 I__2251 (
            .O(N__9101),
            .I(\uut.m6 ));
    Odrv12 I__2250 (
            .O(N__9098),
            .I(\uut.m6 ));
    Odrv4 I__2249 (
            .O(N__9095),
            .I(\uut.m6 ));
    LocalMux I__2248 (
            .O(N__9092),
            .I(\uut.m6 ));
    CascadeMux I__2247 (
            .O(N__9079),
            .I(N__9068));
    InMux I__2246 (
            .O(N__9078),
            .I(N__9065));
    InMux I__2245 (
            .O(N__9077),
            .I(N__9058));
    InMux I__2244 (
            .O(N__9076),
            .I(N__9058));
    InMux I__2243 (
            .O(N__9075),
            .I(N__9058));
    InMux I__2242 (
            .O(N__9074),
            .I(N__9055));
    InMux I__2241 (
            .O(N__9073),
            .I(N__9050));
    InMux I__2240 (
            .O(N__9072),
            .I(N__9047));
    CascadeMux I__2239 (
            .O(N__9071),
            .I(N__9039));
    InMux I__2238 (
            .O(N__9068),
            .I(N__9034));
    LocalMux I__2237 (
            .O(N__9065),
            .I(N__9029));
    LocalMux I__2236 (
            .O(N__9058),
            .I(N__9026));
    LocalMux I__2235 (
            .O(N__9055),
            .I(N__9023));
    InMux I__2234 (
            .O(N__9054),
            .I(N__9020));
    InMux I__2233 (
            .O(N__9053),
            .I(N__9017));
    LocalMux I__2232 (
            .O(N__9050),
            .I(N__9012));
    LocalMux I__2231 (
            .O(N__9047),
            .I(N__9012));
    InMux I__2230 (
            .O(N__9046),
            .I(N__9009));
    InMux I__2229 (
            .O(N__9045),
            .I(N__9006));
    InMux I__2228 (
            .O(N__9044),
            .I(N__9002));
    InMux I__2227 (
            .O(N__9043),
            .I(N__8995));
    InMux I__2226 (
            .O(N__9042),
            .I(N__8995));
    InMux I__2225 (
            .O(N__9039),
            .I(N__8995));
    InMux I__2224 (
            .O(N__9038),
            .I(N__8992));
    InMux I__2223 (
            .O(N__9037),
            .I(N__8989));
    LocalMux I__2222 (
            .O(N__9034),
            .I(N__8986));
    InMux I__2221 (
            .O(N__9033),
            .I(N__8981));
    InMux I__2220 (
            .O(N__9032),
            .I(N__8978));
    Span4Mux_h I__2219 (
            .O(N__9029),
            .I(N__8968));
    Span4Mux_v I__2218 (
            .O(N__9026),
            .I(N__8961));
    Span4Mux_v I__2217 (
            .O(N__9023),
            .I(N__8961));
    LocalMux I__2216 (
            .O(N__9020),
            .I(N__8961));
    LocalMux I__2215 (
            .O(N__9017),
            .I(N__8954));
    Span4Mux_v I__2214 (
            .O(N__9012),
            .I(N__8954));
    LocalMux I__2213 (
            .O(N__9009),
            .I(N__8954));
    LocalMux I__2212 (
            .O(N__9006),
            .I(N__8951));
    InMux I__2211 (
            .O(N__9005),
            .I(N__8948));
    LocalMux I__2210 (
            .O(N__9002),
            .I(N__8941));
    LocalMux I__2209 (
            .O(N__8995),
            .I(N__8941));
    LocalMux I__2208 (
            .O(N__8992),
            .I(N__8941));
    LocalMux I__2207 (
            .O(N__8989),
            .I(N__8938));
    Span4Mux_v I__2206 (
            .O(N__8986),
            .I(N__8935));
    InMux I__2205 (
            .O(N__8985),
            .I(N__8932));
    InMux I__2204 (
            .O(N__8984),
            .I(N__8929));
    LocalMux I__2203 (
            .O(N__8981),
            .I(N__8924));
    LocalMux I__2202 (
            .O(N__8978),
            .I(N__8924));
    InMux I__2201 (
            .O(N__8977),
            .I(N__8920));
    InMux I__2200 (
            .O(N__8976),
            .I(N__8917));
    InMux I__2199 (
            .O(N__8975),
            .I(N__8908));
    InMux I__2198 (
            .O(N__8974),
            .I(N__8908));
    InMux I__2197 (
            .O(N__8973),
            .I(N__8908));
    InMux I__2196 (
            .O(N__8972),
            .I(N__8908));
    InMux I__2195 (
            .O(N__8971),
            .I(N__8905));
    Sp12to4 I__2194 (
            .O(N__8968),
            .I(N__8902));
    Span4Mux_h I__2193 (
            .O(N__8961),
            .I(N__8897));
    Span4Mux_h I__2192 (
            .O(N__8954),
            .I(N__8897));
    Span12Mux_v I__2191 (
            .O(N__8951),
            .I(N__8892));
    LocalMux I__2190 (
            .O(N__8948),
            .I(N__8892));
    Span12Mux_s10_h I__2189 (
            .O(N__8941),
            .I(N__8889));
    Span4Mux_h I__2188 (
            .O(N__8938),
            .I(N__8880));
    Span4Mux_h I__2187 (
            .O(N__8935),
            .I(N__8880));
    LocalMux I__2186 (
            .O(N__8932),
            .I(N__8880));
    LocalMux I__2185 (
            .O(N__8929),
            .I(N__8880));
    Span4Mux_s1_h I__2184 (
            .O(N__8924),
            .I(N__8877));
    InMux I__2183 (
            .O(N__8923),
            .I(N__8874));
    LocalMux I__2182 (
            .O(N__8920),
            .I(\uut.ROM_OE ));
    LocalMux I__2181 (
            .O(N__8917),
            .I(\uut.ROM_OE ));
    LocalMux I__2180 (
            .O(N__8908),
            .I(\uut.ROM_OE ));
    LocalMux I__2179 (
            .O(N__8905),
            .I(\uut.ROM_OE ));
    Odrv12 I__2178 (
            .O(N__8902),
            .I(\uut.ROM_OE ));
    Odrv4 I__2177 (
            .O(N__8897),
            .I(\uut.ROM_OE ));
    Odrv12 I__2176 (
            .O(N__8892),
            .I(\uut.ROM_OE ));
    Odrv12 I__2175 (
            .O(N__8889),
            .I(\uut.ROM_OE ));
    Odrv4 I__2174 (
            .O(N__8880),
            .I(\uut.ROM_OE ));
    Odrv4 I__2173 (
            .O(N__8877),
            .I(\uut.ROM_OE ));
    LocalMux I__2172 (
            .O(N__8874),
            .I(\uut.ROM_OE ));
    InMux I__2171 (
            .O(N__8851),
            .I(N__8833));
    InMux I__2170 (
            .O(N__8850),
            .I(N__8833));
    InMux I__2169 (
            .O(N__8849),
            .I(N__8833));
    InMux I__2168 (
            .O(N__8848),
            .I(N__8833));
    InMux I__2167 (
            .O(N__8847),
            .I(N__8828));
    InMux I__2166 (
            .O(N__8846),
            .I(N__8828));
    InMux I__2165 (
            .O(N__8845),
            .I(N__8822));
    InMux I__2164 (
            .O(N__8844),
            .I(N__8822));
    InMux I__2163 (
            .O(N__8843),
            .I(N__8817));
    InMux I__2162 (
            .O(N__8842),
            .I(N__8817));
    LocalMux I__2161 (
            .O(N__8833),
            .I(N__8812));
    LocalMux I__2160 (
            .O(N__8828),
            .I(N__8812));
    InMux I__2159 (
            .O(N__8827),
            .I(N__8809));
    LocalMux I__2158 (
            .O(N__8822),
            .I(\uut.mar_out_0 ));
    LocalMux I__2157 (
            .O(N__8817),
            .I(\uut.mar_out_0 ));
    Odrv4 I__2156 (
            .O(N__8812),
            .I(\uut.mar_out_0 ));
    LocalMux I__2155 (
            .O(N__8809),
            .I(\uut.mar_out_0 ));
    CEMux I__2154 (
            .O(N__8800),
            .I(N__8796));
    CEMux I__2153 (
            .O(N__8799),
            .I(N__8793));
    LocalMux I__2152 (
            .O(N__8796),
            .I(N__8790));
    LocalMux I__2151 (
            .O(N__8793),
            .I(N__8787));
    Span4Mux_v I__2150 (
            .O(N__8790),
            .I(N__8784));
    Span4Mux_v I__2149 (
            .O(N__8787),
            .I(N__8781));
    Span4Mux_s0_v I__2148 (
            .O(N__8784),
            .I(N__8778));
    Odrv4 I__2147 (
            .O(N__8781),
            .I(\uut.mar.MAR_LD_0_1 ));
    Odrv4 I__2146 (
            .O(N__8778),
            .I(\uut.mar.MAR_LD_0_1 ));
    CascadeMux I__2145 (
            .O(N__8773),
            .I(N__8770));
    InMux I__2144 (
            .O(N__8770),
            .I(N__8762));
    CascadeMux I__2143 (
            .O(N__8769),
            .I(N__8758));
    InMux I__2142 (
            .O(N__8768),
            .I(N__8753));
    InMux I__2141 (
            .O(N__8767),
            .I(N__8750));
    InMux I__2140 (
            .O(N__8766),
            .I(N__8745));
    InMux I__2139 (
            .O(N__8765),
            .I(N__8745));
    LocalMux I__2138 (
            .O(N__8762),
            .I(N__8741));
    InMux I__2137 (
            .O(N__8761),
            .I(N__8736));
    InMux I__2136 (
            .O(N__8758),
            .I(N__8736));
    InMux I__2135 (
            .O(N__8757),
            .I(N__8733));
    InMux I__2134 (
            .O(N__8756),
            .I(N__8730));
    LocalMux I__2133 (
            .O(N__8753),
            .I(N__8727));
    LocalMux I__2132 (
            .O(N__8750),
            .I(N__8724));
    LocalMux I__2131 (
            .O(N__8745),
            .I(N__8721));
    InMux I__2130 (
            .O(N__8744),
            .I(N__8718));
    Span4Mux_h I__2129 (
            .O(N__8741),
            .I(N__8710));
    LocalMux I__2128 (
            .O(N__8736),
            .I(N__8710));
    LocalMux I__2127 (
            .O(N__8733),
            .I(N__8707));
    LocalMux I__2126 (
            .O(N__8730),
            .I(N__8704));
    Span4Mux_v I__2125 (
            .O(N__8727),
            .I(N__8695));
    Span4Mux_v I__2124 (
            .O(N__8724),
            .I(N__8695));
    Span4Mux_s0_h I__2123 (
            .O(N__8721),
            .I(N__8695));
    LocalMux I__2122 (
            .O(N__8718),
            .I(N__8695));
    CascadeMux I__2121 (
            .O(N__8717),
            .I(N__8692));
    CascadeMux I__2120 (
            .O(N__8716),
            .I(N__8689));
    InMux I__2119 (
            .O(N__8715),
            .I(N__8686));
    Span4Mux_v I__2118 (
            .O(N__8710),
            .I(N__8683));
    Span4Mux_v I__2117 (
            .O(N__8707),
            .I(N__8676));
    Span4Mux_v I__2116 (
            .O(N__8704),
            .I(N__8676));
    Span4Mux_h I__2115 (
            .O(N__8695),
            .I(N__8676));
    InMux I__2114 (
            .O(N__8692),
            .I(N__8673));
    InMux I__2113 (
            .O(N__8689),
            .I(N__8670));
    LocalMux I__2112 (
            .O(N__8686),
            .I(\uut.T_2 ));
    Odrv4 I__2111 (
            .O(N__8683),
            .I(\uut.T_2 ));
    Odrv4 I__2110 (
            .O(N__8676),
            .I(\uut.T_2 ));
    LocalMux I__2109 (
            .O(N__8673),
            .I(\uut.T_2 ));
    LocalMux I__2108 (
            .O(N__8670),
            .I(\uut.T_2 ));
    InMux I__2107 (
            .O(N__8659),
            .I(N__8651));
    InMux I__2106 (
            .O(N__8658),
            .I(N__8648));
    InMux I__2105 (
            .O(N__8657),
            .I(N__8643));
    InMux I__2104 (
            .O(N__8656),
            .I(N__8643));
    InMux I__2103 (
            .O(N__8655),
            .I(N__8638));
    InMux I__2102 (
            .O(N__8654),
            .I(N__8638));
    LocalMux I__2101 (
            .O(N__8651),
            .I(N__8635));
    LocalMux I__2100 (
            .O(N__8648),
            .I(N__8630));
    LocalMux I__2099 (
            .O(N__8643),
            .I(N__8627));
    LocalMux I__2098 (
            .O(N__8638),
            .I(N__8624));
    Span12Mux_s11_h I__2097 (
            .O(N__8635),
            .I(N__8621));
    InMux I__2096 (
            .O(N__8634),
            .I(N__8616));
    InMux I__2095 (
            .O(N__8633),
            .I(N__8616));
    Span4Mux_v I__2094 (
            .O(N__8630),
            .I(N__8611));
    Span4Mux_v I__2093 (
            .O(N__8627),
            .I(N__8611));
    Odrv4 I__2092 (
            .O(N__8624),
            .I(\uut.T_0 ));
    Odrv12 I__2091 (
            .O(N__8621),
            .I(\uut.T_0 ));
    LocalMux I__2090 (
            .O(N__8616),
            .I(\uut.T_0 ));
    Odrv4 I__2089 (
            .O(N__8611),
            .I(\uut.T_0 ));
    InMux I__2088 (
            .O(N__8602),
            .I(N__8598));
    CascadeMux I__2087 (
            .O(N__8601),
            .I(N__8594));
    LocalMux I__2086 (
            .O(N__8598),
            .I(N__8591));
    InMux I__2085 (
            .O(N__8597),
            .I(N__8586));
    InMux I__2084 (
            .O(N__8594),
            .I(N__8586));
    Odrv4 I__2083 (
            .O(N__8591),
            .I(\uut.program_counter_3 ));
    LocalMux I__2082 (
            .O(N__8586),
            .I(\uut.program_counter_3 ));
    InMux I__2081 (
            .O(N__8581),
            .I(N__8569));
    InMux I__2080 (
            .O(N__8580),
            .I(N__8569));
    InMux I__2079 (
            .O(N__8579),
            .I(N__8566));
    InMux I__2078 (
            .O(N__8578),
            .I(N__8559));
    InMux I__2077 (
            .O(N__8577),
            .I(N__8559));
    InMux I__2076 (
            .O(N__8576),
            .I(N__8559));
    InMux I__2075 (
            .O(N__8575),
            .I(N__8556));
    InMux I__2074 (
            .O(N__8574),
            .I(N__8553));
    LocalMux I__2073 (
            .O(N__8569),
            .I(N__8546));
    LocalMux I__2072 (
            .O(N__8566),
            .I(N__8541));
    LocalMux I__2071 (
            .O(N__8559),
            .I(N__8541));
    LocalMux I__2070 (
            .O(N__8556),
            .I(N__8536));
    LocalMux I__2069 (
            .O(N__8553),
            .I(N__8536));
    InMux I__2068 (
            .O(N__8552),
            .I(N__8531));
    InMux I__2067 (
            .O(N__8551),
            .I(N__8531));
    InMux I__2066 (
            .O(N__8550),
            .I(N__8528));
    InMux I__2065 (
            .O(N__8549),
            .I(N__8525));
    Span4Mux_v I__2064 (
            .O(N__8546),
            .I(N__8522));
    Span4Mux_h I__2063 (
            .O(N__8541),
            .I(N__8515));
    Span4Mux_s3_h I__2062 (
            .O(N__8536),
            .I(N__8515));
    LocalMux I__2061 (
            .O(N__8531),
            .I(N__8515));
    LocalMux I__2060 (
            .O(N__8528),
            .I(N__8510));
    LocalMux I__2059 (
            .O(N__8525),
            .I(N__8510));
    Odrv4 I__2058 (
            .O(N__8522),
            .I(\uut.D_6 ));
    Odrv4 I__2057 (
            .O(N__8515),
            .I(\uut.D_6 ));
    Odrv12 I__2056 (
            .O(N__8510),
            .I(\uut.D_6 ));
    InMux I__2055 (
            .O(N__8503),
            .I(N__8500));
    LocalMux I__2054 (
            .O(N__8500),
            .I(\uut.program_counter_m_3 ));
    CascadeMux I__2053 (
            .O(N__8497),
            .I(N__8492));
    CascadeMux I__2052 (
            .O(N__8496),
            .I(N__8489));
    InMux I__2051 (
            .O(N__8495),
            .I(N__8485));
    InMux I__2050 (
            .O(N__8492),
            .I(N__8482));
    InMux I__2049 (
            .O(N__8489),
            .I(N__8479));
    InMux I__2048 (
            .O(N__8488),
            .I(N__8474));
    LocalMux I__2047 (
            .O(N__8485),
            .I(N__8471));
    LocalMux I__2046 (
            .O(N__8482),
            .I(N__8466));
    LocalMux I__2045 (
            .O(N__8479),
            .I(N__8466));
    CascadeMux I__2044 (
            .O(N__8478),
            .I(N__8461));
    InMux I__2043 (
            .O(N__8477),
            .I(N__8458));
    LocalMux I__2042 (
            .O(N__8474),
            .I(N__8455));
    Span4Mux_h I__2041 (
            .O(N__8471),
            .I(N__8450));
    Span4Mux_v I__2040 (
            .O(N__8466),
            .I(N__8450));
    InMux I__2039 (
            .O(N__8465),
            .I(N__8445));
    InMux I__2038 (
            .O(N__8464),
            .I(N__8445));
    InMux I__2037 (
            .O(N__8461),
            .I(N__8442));
    LocalMux I__2036 (
            .O(N__8458),
            .I(\uut.acc_out_3 ));
    Odrv12 I__2035 (
            .O(N__8455),
            .I(\uut.acc_out_3 ));
    Odrv4 I__2034 (
            .O(N__8450),
            .I(\uut.acc_out_3 ));
    LocalMux I__2033 (
            .O(N__8445),
            .I(\uut.acc_out_3 ));
    LocalMux I__2032 (
            .O(N__8442),
            .I(\uut.acc_out_3 ));
    CascadeMux I__2031 (
            .O(N__8431),
            .I(N__8427));
    InMux I__2030 (
            .O(N__8430),
            .I(N__8423));
    InMux I__2029 (
            .O(N__8427),
            .I(N__8420));
    InMux I__2028 (
            .O(N__8426),
            .I(N__8417));
    LocalMux I__2027 (
            .O(N__8423),
            .I(N__8411));
    LocalMux I__2026 (
            .O(N__8420),
            .I(N__8411));
    LocalMux I__2025 (
            .O(N__8417),
            .I(N__8408));
    CascadeMux I__2024 (
            .O(N__8416),
            .I(N__8405));
    Span4Mux_v I__2023 (
            .O(N__8411),
            .I(N__8401));
    Span4Mux_s3_h I__2022 (
            .O(N__8408),
            .I(N__8398));
    InMux I__2021 (
            .O(N__8405),
            .I(N__8393));
    InMux I__2020 (
            .O(N__8404),
            .I(N__8393));
    Odrv4 I__2019 (
            .O(N__8401),
            .I(\uut.ir_out_3 ));
    Odrv4 I__2018 (
            .O(N__8398),
            .I(\uut.ir_out_3 ));
    LocalMux I__2017 (
            .O(N__8393),
            .I(\uut.ir_out_3 ));
    InMux I__2016 (
            .O(N__8386),
            .I(N__8379));
    InMux I__2015 (
            .O(N__8385),
            .I(N__8376));
    InMux I__2014 (
            .O(N__8384),
            .I(N__8372));
    InMux I__2013 (
            .O(N__8383),
            .I(N__8369));
    InMux I__2012 (
            .O(N__8382),
            .I(N__8366));
    LocalMux I__2011 (
            .O(N__8379),
            .I(N__8361));
    LocalMux I__2010 (
            .O(N__8376),
            .I(N__8361));
    InMux I__2009 (
            .O(N__8375),
            .I(N__8356));
    LocalMux I__2008 (
            .O(N__8372),
            .I(N__8353));
    LocalMux I__2007 (
            .O(N__8369),
            .I(N__8350));
    LocalMux I__2006 (
            .O(N__8366),
            .I(N__8347));
    Span4Mux_h I__2005 (
            .O(N__8361),
            .I(N__8344));
    InMux I__2004 (
            .O(N__8360),
            .I(N__8341));
    InMux I__2003 (
            .O(N__8359),
            .I(N__8338));
    LocalMux I__2002 (
            .O(N__8356),
            .I(N__8335));
    Span4Mux_s2_h I__2001 (
            .O(N__8353),
            .I(N__8332));
    Span4Mux_s2_h I__2000 (
            .O(N__8350),
            .I(N__8329));
    Span4Mux_s3_h I__1999 (
            .O(N__8347),
            .I(N__8324));
    Span4Mux_v I__1998 (
            .O(N__8344),
            .I(N__8324));
    LocalMux I__1997 (
            .O(N__8341),
            .I(N__8321));
    LocalMux I__1996 (
            .O(N__8338),
            .I(\uut.un5_MAR_LD ));
    Odrv4 I__1995 (
            .O(N__8335),
            .I(\uut.un5_MAR_LD ));
    Odrv4 I__1994 (
            .O(N__8332),
            .I(\uut.un5_MAR_LD ));
    Odrv4 I__1993 (
            .O(N__8329),
            .I(\uut.un5_MAR_LD ));
    Odrv4 I__1992 (
            .O(N__8324),
            .I(\uut.un5_MAR_LD ));
    Odrv12 I__1991 (
            .O(N__8321),
            .I(\uut.un5_MAR_LD ));
    CascadeMux I__1990 (
            .O(N__8308),
            .I(\uut.AR_BUF.out_1_ivZ0Z_0_cascade_ ));
    InMux I__1989 (
            .O(N__8305),
            .I(N__8302));
    LocalMux I__1988 (
            .O(N__8302),
            .I(N__8298));
    InMux I__1987 (
            .O(N__8301),
            .I(N__8295));
    Odrv4 I__1986 (
            .O(N__8298),
            .I(\uut.out_1_iv_2 ));
    LocalMux I__1985 (
            .O(N__8295),
            .I(\uut.out_1_iv_2 ));
    CascadeMux I__1984 (
            .O(N__8290),
            .I(\uut.out_1_iv_2_1_cascade_ ));
    InMux I__1983 (
            .O(N__8287),
            .I(N__8283));
    InMux I__1982 (
            .O(N__8286),
            .I(N__8275));
    LocalMux I__1981 (
            .O(N__8283),
            .I(N__8268));
    InMux I__1980 (
            .O(N__8282),
            .I(N__8265));
    InMux I__1979 (
            .O(N__8281),
            .I(N__8262));
    InMux I__1978 (
            .O(N__8280),
            .I(N__8257));
    InMux I__1977 (
            .O(N__8279),
            .I(N__8254));
    InMux I__1976 (
            .O(N__8278),
            .I(N__8250));
    LocalMux I__1975 (
            .O(N__8275),
            .I(N__8247));
    InMux I__1974 (
            .O(N__8274),
            .I(N__8242));
    InMux I__1973 (
            .O(N__8273),
            .I(N__8242));
    InMux I__1972 (
            .O(N__8272),
            .I(N__8239));
    InMux I__1971 (
            .O(N__8271),
            .I(N__8236));
    Span4Mux_h I__1970 (
            .O(N__8268),
            .I(N__8229));
    LocalMux I__1969 (
            .O(N__8265),
            .I(N__8229));
    LocalMux I__1968 (
            .O(N__8262),
            .I(N__8229));
    InMux I__1967 (
            .O(N__8261),
            .I(N__8226));
    InMux I__1966 (
            .O(N__8260),
            .I(N__8223));
    LocalMux I__1965 (
            .O(N__8257),
            .I(N__8218));
    LocalMux I__1964 (
            .O(N__8254),
            .I(N__8218));
    InMux I__1963 (
            .O(N__8253),
            .I(N__8215));
    LocalMux I__1962 (
            .O(N__8250),
            .I(N__8210));
    Span4Mux_v I__1961 (
            .O(N__8247),
            .I(N__8210));
    LocalMux I__1960 (
            .O(N__8242),
            .I(N__8205));
    LocalMux I__1959 (
            .O(N__8239),
            .I(N__8205));
    LocalMux I__1958 (
            .O(N__8236),
            .I(N__8200));
    Span4Mux_v I__1957 (
            .O(N__8229),
            .I(N__8200));
    LocalMux I__1956 (
            .O(N__8226),
            .I(N__8197));
    LocalMux I__1955 (
            .O(N__8223),
            .I(N__8194));
    Span4Mux_v I__1954 (
            .O(N__8218),
            .I(N__8191));
    LocalMux I__1953 (
            .O(N__8215),
            .I(N__8188));
    Span4Mux_v I__1952 (
            .O(N__8210),
            .I(N__8183));
    Span4Mux_h I__1951 (
            .O(N__8205),
            .I(N__8183));
    Span4Mux_h I__1950 (
            .O(N__8200),
            .I(N__8178));
    Span4Mux_s2_h I__1949 (
            .O(N__8197),
            .I(N__8178));
    Span12Mux_s8_h I__1948 (
            .O(N__8194),
            .I(N__8175));
    Sp12to4 I__1947 (
            .O(N__8191),
            .I(N__8170));
    Span12Mux_v I__1946 (
            .O(N__8188),
            .I(N__8170));
    Odrv4 I__1945 (
            .O(N__8183),
            .I(\uut.OUT_LD ));
    Odrv4 I__1944 (
            .O(N__8178),
            .I(\uut.OUT_LD ));
    Odrv12 I__1943 (
            .O(N__8175),
            .I(\uut.OUT_LD ));
    Odrv12 I__1942 (
            .O(N__8170),
            .I(\uut.OUT_LD ));
    IoInMux I__1941 (
            .O(N__8161),
            .I(N__8158));
    LocalMux I__1940 (
            .O(N__8158),
            .I(N__8154));
    InMux I__1939 (
            .O(N__8157),
            .I(N__8151));
    Span12Mux_s0_h I__1938 (
            .O(N__8154),
            .I(N__8148));
    LocalMux I__1937 (
            .O(N__8151),
            .I(N__8145));
    Odrv12 I__1936 (
            .O(N__8148),
            .I(LED4_c));
    Odrv4 I__1935 (
            .O(N__8145),
            .I(LED4_c));
    InMux I__1934 (
            .O(N__8140),
            .I(N__8137));
    LocalMux I__1933 (
            .O(N__8137),
            .I(\uut.alu_out_m_3 ));
    CascadeMux I__1932 (
            .O(N__8134),
            .I(\uut.m15_cascade_ ));
    InMux I__1931 (
            .O(N__8131),
            .I(N__8128));
    LocalMux I__1930 (
            .O(N__8128),
            .I(\uut.out_1_iv_3 ));
    CascadeMux I__1929 (
            .O(N__8125),
            .I(N__8122));
    InMux I__1928 (
            .O(N__8122),
            .I(N__8118));
    InMux I__1927 (
            .O(N__8121),
            .I(N__8115));
    LocalMux I__1926 (
            .O(N__8118),
            .I(N__8112));
    LocalMux I__1925 (
            .O(N__8115),
            .I(N__8109));
    Span4Mux_s3_v I__1924 (
            .O(N__8112),
            .I(N__8103));
    Span4Mux_s0_h I__1923 (
            .O(N__8109),
            .I(N__8103));
    InMux I__1922 (
            .O(N__8108),
            .I(N__8100));
    Span4Mux_h I__1921 (
            .O(N__8103),
            .I(N__8095));
    LocalMux I__1920 (
            .O(N__8100),
            .I(N__8092));
    InMux I__1919 (
            .O(N__8099),
            .I(N__8089));
    InMux I__1918 (
            .O(N__8098),
            .I(N__8086));
    Odrv4 I__1917 (
            .O(N__8095),
            .I(\uut.out_1_0_ivdup_2 ));
    Odrv12 I__1916 (
            .O(N__8092),
            .I(\uut.out_1_0_ivdup_2 ));
    LocalMux I__1915 (
            .O(N__8089),
            .I(\uut.out_1_0_ivdup_2 ));
    LocalMux I__1914 (
            .O(N__8086),
            .I(\uut.out_1_0_ivdup_2 ));
    InMux I__1913 (
            .O(N__8077),
            .I(N__8074));
    LocalMux I__1912 (
            .O(N__8074),
            .I(N__8070));
    InMux I__1911 (
            .O(N__8073),
            .I(N__8067));
    Span4Mux_s3_v I__1910 (
            .O(N__8070),
            .I(N__8063));
    LocalMux I__1909 (
            .O(N__8067),
            .I(N__8060));
    InMux I__1908 (
            .O(N__8066),
            .I(N__8057));
    Span4Mux_h I__1907 (
            .O(N__8063),
            .I(N__8050));
    Span4Mux_s3_v I__1906 (
            .O(N__8060),
            .I(N__8050));
    LocalMux I__1905 (
            .O(N__8057),
            .I(N__8050));
    Odrv4 I__1904 (
            .O(N__8050),
            .I(\uut.out_1_0_iv_3 ));
    CascadeMux I__1903 (
            .O(N__8047),
            .I(N__8044));
    InMux I__1902 (
            .O(N__8044),
            .I(N__8038));
    InMux I__1901 (
            .O(N__8043),
            .I(N__8038));
    LocalMux I__1900 (
            .O(N__8038),
            .I(N__8035));
    Odrv12 I__1899 (
            .O(N__8035),
            .I(\uut.MAR_LD_0 ));
    InMux I__1898 (
            .O(N__8032),
            .I(N__8028));
    CEMux I__1897 (
            .O(N__8031),
            .I(N__8024));
    LocalMux I__1896 (
            .O(N__8028),
            .I(N__8020));
    CEMux I__1895 (
            .O(N__8027),
            .I(N__8017));
    LocalMux I__1894 (
            .O(N__8024),
            .I(N__8014));
    InMux I__1893 (
            .O(N__8023),
            .I(N__8011));
    Span4Mux_h I__1892 (
            .O(N__8020),
            .I(N__8008));
    LocalMux I__1891 (
            .O(N__8017),
            .I(N__8005));
    Span4Mux_s0_h I__1890 (
            .O(N__8014),
            .I(N__8002));
    LocalMux I__1889 (
            .O(N__8011),
            .I(N__7999));
    Span4Mux_h I__1888 (
            .O(N__8008),
            .I(N__7996));
    Odrv12 I__1887 (
            .O(N__8005),
            .I(\uut.AR_LD ));
    Odrv4 I__1886 (
            .O(N__8002),
            .I(\uut.AR_LD ));
    Odrv4 I__1885 (
            .O(N__7999),
            .I(\uut.AR_LD ));
    Odrv4 I__1884 (
            .O(N__7996),
            .I(\uut.AR_LD ));
    InMux I__1883 (
            .O(N__7987),
            .I(N__7982));
    InMux I__1882 (
            .O(N__7986),
            .I(N__7979));
    InMux I__1881 (
            .O(N__7985),
            .I(N__7976));
    LocalMux I__1880 (
            .O(N__7982),
            .I(N__7971));
    LocalMux I__1879 (
            .O(N__7979),
            .I(N__7966));
    LocalMux I__1878 (
            .O(N__7976),
            .I(N__7966));
    CascadeMux I__1877 (
            .O(N__7975),
            .I(N__7962));
    InMux I__1876 (
            .O(N__7974),
            .I(N__7959));
    Span4Mux_v I__1875 (
            .O(N__7971),
            .I(N__7954));
    Span4Mux_v I__1874 (
            .O(N__7966),
            .I(N__7954));
    InMux I__1873 (
            .O(N__7965),
            .I(N__7949));
    InMux I__1872 (
            .O(N__7962),
            .I(N__7949));
    LocalMux I__1871 (
            .O(N__7959),
            .I(N__7946));
    Odrv4 I__1870 (
            .O(N__7954),
            .I(\uut.un14_MAR_LD ));
    LocalMux I__1869 (
            .O(N__7949),
            .I(\uut.un14_MAR_LD ));
    Odrv4 I__1868 (
            .O(N__7946),
            .I(\uut.un14_MAR_LD ));
    InMux I__1867 (
            .O(N__7939),
            .I(N__7936));
    LocalMux I__1866 (
            .O(N__7936),
            .I(N__7930));
    InMux I__1865 (
            .O(N__7935),
            .I(N__7926));
    InMux I__1864 (
            .O(N__7934),
            .I(N__7921));
    InMux I__1863 (
            .O(N__7933),
            .I(N__7921));
    Span4Mux_s1_h I__1862 (
            .O(N__7930),
            .I(N__7918));
    InMux I__1861 (
            .O(N__7929),
            .I(N__7915));
    LocalMux I__1860 (
            .O(N__7926),
            .I(N__7912));
    LocalMux I__1859 (
            .O(N__7921),
            .I(N__7909));
    Span4Mux_v I__1858 (
            .O(N__7918),
            .I(N__7904));
    LocalMux I__1857 (
            .O(N__7915),
            .I(N__7904));
    Span4Mux_s3_h I__1856 (
            .O(N__7912),
            .I(N__7899));
    Span4Mux_h I__1855 (
            .O(N__7909),
            .I(N__7899));
    Odrv4 I__1854 (
            .O(N__7904),
            .I(\uut.un8_MAR_LD ));
    Odrv4 I__1853 (
            .O(N__7899),
            .I(\uut.un8_MAR_LD ));
    InMux I__1852 (
            .O(N__7894),
            .I(N__7889));
    InMux I__1851 (
            .O(N__7893),
            .I(N__7886));
    InMux I__1850 (
            .O(N__7892),
            .I(N__7883));
    LocalMux I__1849 (
            .O(N__7889),
            .I(N__7880));
    LocalMux I__1848 (
            .O(N__7886),
            .I(N__7877));
    LocalMux I__1847 (
            .O(N__7883),
            .I(N__7874));
    Span4Mux_s3_v I__1846 (
            .O(N__7880),
            .I(N__7869));
    Span4Mux_v I__1845 (
            .O(N__7877),
            .I(N__7864));
    Span4Mux_s3_h I__1844 (
            .O(N__7874),
            .I(N__7864));
    InMux I__1843 (
            .O(N__7873),
            .I(N__7859));
    InMux I__1842 (
            .O(N__7872),
            .I(N__7859));
    Odrv4 I__1841 (
            .O(N__7869),
            .I(\uut.un1_IR_OE_4_1 ));
    Odrv4 I__1840 (
            .O(N__7864),
            .I(\uut.un1_IR_OE_4_1 ));
    LocalMux I__1839 (
            .O(N__7859),
            .I(\uut.un1_IR_OE_4_1 ));
    InMux I__1838 (
            .O(N__7852),
            .I(N__7849));
    LocalMux I__1837 (
            .O(N__7849),
            .I(\uut.pc.un1_inc_0_0 ));
    CascadeMux I__1836 (
            .O(N__7846),
            .I(\uut.ir_out_m_d_3_cascade_ ));
    InMux I__1835 (
            .O(N__7843),
            .I(N__7840));
    LocalMux I__1834 (
            .O(N__7840),
            .I(\uut.pc.g0_sn ));
    InMux I__1833 (
            .O(N__7837),
            .I(N__7833));
    InMux I__1832 (
            .O(N__7836),
            .I(N__7830));
    LocalMux I__1831 (
            .O(N__7833),
            .I(N__7827));
    LocalMux I__1830 (
            .O(N__7830),
            .I(N__7824));
    Span12Mux_s10_h I__1829 (
            .O(N__7827),
            .I(N__7821));
    Span4Mux_v I__1828 (
            .O(N__7824),
            .I(N__7818));
    Odrv12 I__1827 (
            .O(N__7821),
            .I(\uut.seq.counter.T_1Z0Z_4 ));
    Odrv4 I__1826 (
            .O(N__7818),
            .I(\uut.seq.counter.T_1Z0Z_4 ));
    CascadeMux I__1825 (
            .O(N__7813),
            .I(\uut.AR_BUF.out_1_ivdupZ0Z_0_cascade_ ));
    InMux I__1824 (
            .O(N__7810),
            .I(N__7807));
    LocalMux I__1823 (
            .O(N__7807),
            .I(\uut.g0_0 ));
    InMux I__1822 (
            .O(N__7804),
            .I(N__7800));
    CascadeMux I__1821 (
            .O(N__7803),
            .I(N__7797));
    LocalMux I__1820 (
            .O(N__7800),
            .I(N__7794));
    InMux I__1819 (
            .O(N__7797),
            .I(N__7791));
    Odrv4 I__1818 (
            .O(N__7794),
            .I(\uut.AR_out_3 ));
    LocalMux I__1817 (
            .O(N__7791),
            .I(\uut.AR_out_3 ));
    CascadeMux I__1816 (
            .O(N__7786),
            .I(\uut.g1_cascade_ ));
    InMux I__1815 (
            .O(N__7783),
            .I(N__7776));
    InMux I__1814 (
            .O(N__7782),
            .I(N__7773));
    InMux I__1813 (
            .O(N__7781),
            .I(N__7770));
    InMux I__1812 (
            .O(N__7780),
            .I(N__7765));
    InMux I__1811 (
            .O(N__7779),
            .I(N__7765));
    LocalMux I__1810 (
            .O(N__7776),
            .I(N__7755));
    LocalMux I__1809 (
            .O(N__7773),
            .I(N__7748));
    LocalMux I__1808 (
            .O(N__7770),
            .I(N__7748));
    LocalMux I__1807 (
            .O(N__7765),
            .I(N__7748));
    InMux I__1806 (
            .O(N__7764),
            .I(N__7745));
    InMux I__1805 (
            .O(N__7763),
            .I(N__7742));
    InMux I__1804 (
            .O(N__7762),
            .I(N__7739));
    InMux I__1803 (
            .O(N__7761),
            .I(N__7736));
    InMux I__1802 (
            .O(N__7760),
            .I(N__7733));
    InMux I__1801 (
            .O(N__7759),
            .I(N__7728));
    InMux I__1800 (
            .O(N__7758),
            .I(N__7728));
    Span4Mux_v I__1799 (
            .O(N__7755),
            .I(N__7725));
    Span4Mux_v I__1798 (
            .O(N__7748),
            .I(N__7722));
    LocalMux I__1797 (
            .O(N__7745),
            .I(N__7715));
    LocalMux I__1796 (
            .O(N__7742),
            .I(N__7715));
    LocalMux I__1795 (
            .O(N__7739),
            .I(N__7715));
    LocalMux I__1794 (
            .O(N__7736),
            .I(N__7708));
    LocalMux I__1793 (
            .O(N__7733),
            .I(N__7708));
    LocalMux I__1792 (
            .O(N__7728),
            .I(N__7708));
    Odrv4 I__1791 (
            .O(N__7725),
            .I(\uut.T_2_rep1_RNI6BLF1 ));
    Odrv4 I__1790 (
            .O(N__7722),
            .I(\uut.T_2_rep1_RNI6BLF1 ));
    Odrv4 I__1789 (
            .O(N__7715),
            .I(\uut.T_2_rep1_RNI6BLF1 ));
    Odrv4 I__1788 (
            .O(N__7708),
            .I(\uut.T_2_rep1_RNI6BLF1 ));
    InMux I__1787 (
            .O(N__7699),
            .I(N__7696));
    LocalMux I__1786 (
            .O(N__7696),
            .I(\uut.AR_BUF.g0_1_0 ));
    InMux I__1785 (
            .O(N__7693),
            .I(N__7689));
    InMux I__1784 (
            .O(N__7692),
            .I(N__7685));
    LocalMux I__1783 (
            .O(N__7689),
            .I(N__7681));
    InMux I__1782 (
            .O(N__7688),
            .I(N__7677));
    LocalMux I__1781 (
            .O(N__7685),
            .I(N__7674));
    InMux I__1780 (
            .O(N__7684),
            .I(N__7671));
    Span4Mux_h I__1779 (
            .O(N__7681),
            .I(N__7668));
    InMux I__1778 (
            .O(N__7680),
            .I(N__7665));
    LocalMux I__1777 (
            .O(N__7677),
            .I(N__7662));
    Span12Mux_s7_v I__1776 (
            .O(N__7674),
            .I(N__7657));
    LocalMux I__1775 (
            .O(N__7671),
            .I(N__7657));
    Span4Mux_v I__1774 (
            .O(N__7668),
            .I(N__7652));
    LocalMux I__1773 (
            .O(N__7665),
            .I(N__7652));
    Odrv12 I__1772 (
            .O(N__7662),
            .I(\uut.alu_out_m_1 ));
    Odrv12 I__1771 (
            .O(N__7657),
            .I(\uut.alu_out_m_1 ));
    Odrv4 I__1770 (
            .O(N__7652),
            .I(\uut.alu_out_m_1 ));
    InMux I__1769 (
            .O(N__7645),
            .I(N__7640));
    InMux I__1768 (
            .O(N__7644),
            .I(N__7637));
    InMux I__1767 (
            .O(N__7643),
            .I(N__7633));
    LocalMux I__1766 (
            .O(N__7640),
            .I(N__7630));
    LocalMux I__1765 (
            .O(N__7637),
            .I(N__7627));
    InMux I__1764 (
            .O(N__7636),
            .I(N__7624));
    LocalMux I__1763 (
            .O(N__7633),
            .I(N__7620));
    Span4Mux_s2_v I__1762 (
            .O(N__7630),
            .I(N__7617));
    Span12Mux_s10_h I__1761 (
            .O(N__7627),
            .I(N__7612));
    LocalMux I__1760 (
            .O(N__7624),
            .I(N__7612));
    InMux I__1759 (
            .O(N__7623),
            .I(N__7609));
    Span12Mux_v I__1758 (
            .O(N__7620),
            .I(N__7606));
    Odrv4 I__1757 (
            .O(N__7617),
            .I(\uut.N_11_i_m ));
    Odrv12 I__1756 (
            .O(N__7612),
            .I(\uut.N_11_i_m ));
    LocalMux I__1755 (
            .O(N__7609),
            .I(\uut.N_11_i_m ));
    Odrv12 I__1754 (
            .O(N__7606),
            .I(\uut.N_11_i_m ));
    InMux I__1753 (
            .O(N__7597),
            .I(N__7593));
    InMux I__1752 (
            .O(N__7596),
            .I(N__7590));
    LocalMux I__1751 (
            .O(N__7593),
            .I(N__7586));
    LocalMux I__1750 (
            .O(N__7590),
            .I(N__7583));
    InMux I__1749 (
            .O(N__7589),
            .I(N__7580));
    Span4Mux_s3_v I__1748 (
            .O(N__7586),
            .I(N__7576));
    Span4Mux_s3_v I__1747 (
            .O(N__7583),
            .I(N__7571));
    LocalMux I__1746 (
            .O(N__7580),
            .I(N__7571));
    InMux I__1745 (
            .O(N__7579),
            .I(N__7568));
    Span4Mux_v I__1744 (
            .O(N__7576),
            .I(N__7562));
    Span4Mux_v I__1743 (
            .O(N__7571),
            .I(N__7562));
    LocalMux I__1742 (
            .O(N__7568),
            .I(N__7559));
    InMux I__1741 (
            .O(N__7567),
            .I(N__7556));
    Odrv4 I__1740 (
            .O(N__7562),
            .I(\uut.out_1_1_iv_3dup_1 ));
    Odrv4 I__1739 (
            .O(N__7559),
            .I(\uut.out_1_1_iv_3dup_1 ));
    LocalMux I__1738 (
            .O(N__7556),
            .I(\uut.out_1_1_iv_3dup_1 ));
    InMux I__1737 (
            .O(N__7549),
            .I(N__7544));
    InMux I__1736 (
            .O(N__7548),
            .I(N__7541));
    InMux I__1735 (
            .O(N__7547),
            .I(N__7538));
    LocalMux I__1734 (
            .O(N__7544),
            .I(N__7535));
    LocalMux I__1733 (
            .O(N__7541),
            .I(N__7532));
    LocalMux I__1732 (
            .O(N__7538),
            .I(N__7529));
    Span4Mux_h I__1731 (
            .O(N__7535),
            .I(N__7526));
    Span4Mux_h I__1730 (
            .O(N__7532),
            .I(N__7523));
    Odrv12 I__1729 (
            .O(N__7529),
            .I(\uut.b_reg_out_1 ));
    Odrv4 I__1728 (
            .O(N__7526),
            .I(\uut.b_reg_out_1 ));
    Odrv4 I__1727 (
            .O(N__7523),
            .I(\uut.b_reg_out_1 ));
    CEMux I__1726 (
            .O(N__7516),
            .I(N__7511));
    CEMux I__1725 (
            .O(N__7515),
            .I(N__7507));
    CEMux I__1724 (
            .O(N__7514),
            .I(N__7504));
    LocalMux I__1723 (
            .O(N__7511),
            .I(N__7500));
    CEMux I__1722 (
            .O(N__7510),
            .I(N__7497));
    LocalMux I__1721 (
            .O(N__7507),
            .I(N__7494));
    LocalMux I__1720 (
            .O(N__7504),
            .I(N__7491));
    CEMux I__1719 (
            .O(N__7503),
            .I(N__7488));
    Span4Mux_h I__1718 (
            .O(N__7500),
            .I(N__7482));
    LocalMux I__1717 (
            .O(N__7497),
            .I(N__7482));
    Span4Mux_v I__1716 (
            .O(N__7494),
            .I(N__7476));
    Span4Mux_v I__1715 (
            .O(N__7491),
            .I(N__7476));
    LocalMux I__1714 (
            .O(N__7488),
            .I(N__7473));
    CEMux I__1713 (
            .O(N__7487),
            .I(N__7470));
    Span4Mux_v I__1712 (
            .O(N__7482),
            .I(N__7467));
    CEMux I__1711 (
            .O(N__7481),
            .I(N__7464));
    Span4Mux_s2_v I__1710 (
            .O(N__7476),
            .I(N__7461));
    Span4Mux_v I__1709 (
            .O(N__7473),
            .I(N__7458));
    LocalMux I__1708 (
            .O(N__7470),
            .I(N__7455));
    Span4Mux_h I__1707 (
            .O(N__7467),
            .I(N__7450));
    LocalMux I__1706 (
            .O(N__7464),
            .I(N__7450));
    Span4Mux_h I__1705 (
            .O(N__7461),
            .I(N__7447));
    Span4Mux_h I__1704 (
            .O(N__7458),
            .I(N__7444));
    Span4Mux_h I__1703 (
            .O(N__7455),
            .I(N__7439));
    Span4Mux_s1_h I__1702 (
            .O(N__7450),
            .I(N__7439));
    Odrv4 I__1701 (
            .O(N__7447),
            .I(\uut.B_LD_0_i ));
    Odrv4 I__1700 (
            .O(N__7444),
            .I(\uut.B_LD_0_i ));
    Odrv4 I__1699 (
            .O(N__7439),
            .I(\uut.B_LD_0_i ));
    CEMux I__1698 (
            .O(N__7432),
            .I(N__7429));
    LocalMux I__1697 (
            .O(N__7429),
            .I(N__7425));
    CEMux I__1696 (
            .O(N__7428),
            .I(N__7422));
    Span4Mux_s2_v I__1695 (
            .O(N__7425),
            .I(N__7407));
    LocalMux I__1694 (
            .O(N__7422),
            .I(N__7407));
    InMux I__1693 (
            .O(N__7421),
            .I(N__7392));
    InMux I__1692 (
            .O(N__7420),
            .I(N__7392));
    InMux I__1691 (
            .O(N__7419),
            .I(N__7392));
    InMux I__1690 (
            .O(N__7418),
            .I(N__7392));
    InMux I__1689 (
            .O(N__7417),
            .I(N__7387));
    InMux I__1688 (
            .O(N__7416),
            .I(N__7387));
    InMux I__1687 (
            .O(N__7415),
            .I(N__7383));
    InMux I__1686 (
            .O(N__7414),
            .I(N__7378));
    InMux I__1685 (
            .O(N__7413),
            .I(N__7378));
    InMux I__1684 (
            .O(N__7412),
            .I(N__7375));
    Span4Mux_v I__1683 (
            .O(N__7407),
            .I(N__7372));
    InMux I__1682 (
            .O(N__7406),
            .I(N__7369));
    InMux I__1681 (
            .O(N__7405),
            .I(N__7364));
    InMux I__1680 (
            .O(N__7404),
            .I(N__7364));
    InMux I__1679 (
            .O(N__7403),
            .I(N__7361));
    InMux I__1678 (
            .O(N__7402),
            .I(N__7357));
    CEMux I__1677 (
            .O(N__7401),
            .I(N__7354));
    LocalMux I__1676 (
            .O(N__7392),
            .I(N__7351));
    LocalMux I__1675 (
            .O(N__7387),
            .I(N__7348));
    InMux I__1674 (
            .O(N__7386),
            .I(N__7345));
    LocalMux I__1673 (
            .O(N__7383),
            .I(N__7340));
    LocalMux I__1672 (
            .O(N__7378),
            .I(N__7340));
    LocalMux I__1671 (
            .O(N__7375),
            .I(N__7329));
    Span4Mux_h I__1670 (
            .O(N__7372),
            .I(N__7329));
    LocalMux I__1669 (
            .O(N__7369),
            .I(N__7329));
    LocalMux I__1668 (
            .O(N__7364),
            .I(N__7329));
    LocalMux I__1667 (
            .O(N__7361),
            .I(N__7329));
    CascadeMux I__1666 (
            .O(N__7360),
            .I(N__7324));
    LocalMux I__1665 (
            .O(N__7357),
            .I(N__7321));
    LocalMux I__1664 (
            .O(N__7354),
            .I(N__7312));
    Span4Mux_s2_v I__1663 (
            .O(N__7351),
            .I(N__7312));
    Span4Mux_s2_v I__1662 (
            .O(N__7348),
            .I(N__7312));
    LocalMux I__1661 (
            .O(N__7345),
            .I(N__7312));
    Span4Mux_v I__1660 (
            .O(N__7340),
            .I(N__7305));
    Span4Mux_v I__1659 (
            .O(N__7329),
            .I(N__7302));
    InMux I__1658 (
            .O(N__7328),
            .I(N__7297));
    InMux I__1657 (
            .O(N__7327),
            .I(N__7297));
    InMux I__1656 (
            .O(N__7324),
            .I(N__7294));
    Span12Mux_s2_v I__1655 (
            .O(N__7321),
            .I(N__7291));
    Span4Mux_v I__1654 (
            .O(N__7312),
            .I(N__7288));
    InMux I__1653 (
            .O(N__7311),
            .I(N__7285));
    InMux I__1652 (
            .O(N__7310),
            .I(N__7278));
    InMux I__1651 (
            .O(N__7309),
            .I(N__7278));
    InMux I__1650 (
            .O(N__7308),
            .I(N__7278));
    Sp12to4 I__1649 (
            .O(N__7305),
            .I(N__7269));
    Sp12to4 I__1648 (
            .O(N__7302),
            .I(N__7269));
    LocalMux I__1647 (
            .O(N__7297),
            .I(N__7269));
    LocalMux I__1646 (
            .O(N__7294),
            .I(N__7269));
    Odrv12 I__1645 (
            .O(N__7291),
            .I(\uut.inc ));
    Odrv4 I__1644 (
            .O(N__7288),
            .I(\uut.inc ));
    LocalMux I__1643 (
            .O(N__7285),
            .I(\uut.inc ));
    LocalMux I__1642 (
            .O(N__7278),
            .I(\uut.inc ));
    Odrv12 I__1641 (
            .O(N__7269),
            .I(\uut.inc ));
    CascadeMux I__1640 (
            .O(N__7258),
            .I(N__7255));
    InMux I__1639 (
            .O(N__7255),
            .I(N__7251));
    CascadeMux I__1638 (
            .O(N__7254),
            .I(N__7248));
    LocalMux I__1637 (
            .O(N__7251),
            .I(N__7244));
    InMux I__1636 (
            .O(N__7248),
            .I(N__7239));
    InMux I__1635 (
            .O(N__7247),
            .I(N__7239));
    Span4Mux_h I__1634 (
            .O(N__7244),
            .I(N__7234));
    LocalMux I__1633 (
            .O(N__7239),
            .I(N__7231));
    InMux I__1632 (
            .O(N__7238),
            .I(N__7228));
    InMux I__1631 (
            .O(N__7237),
            .I(N__7225));
    Span4Mux_v I__1630 (
            .O(N__7234),
            .I(N__7222));
    Span12Mux_v I__1629 (
            .O(N__7231),
            .I(N__7217));
    LocalMux I__1628 (
            .O(N__7228),
            .I(N__7217));
    LocalMux I__1627 (
            .O(N__7225),
            .I(\uut.ir_out_2 ));
    Odrv4 I__1626 (
            .O(N__7222),
            .I(\uut.ir_out_2 ));
    Odrv12 I__1625 (
            .O(N__7217),
            .I(\uut.ir_out_2 ));
    InMux I__1624 (
            .O(N__7210),
            .I(N__7206));
    InMux I__1623 (
            .O(N__7209),
            .I(N__7203));
    LocalMux I__1622 (
            .O(N__7206),
            .I(N__7200));
    LocalMux I__1621 (
            .O(N__7203),
            .I(N__7197));
    Odrv4 I__1620 (
            .O(N__7200),
            .I(\uut.N_14_0 ));
    Odrv4 I__1619 (
            .O(N__7197),
            .I(\uut.N_14_0 ));
    InMux I__1618 (
            .O(N__7192),
            .I(N__7189));
    LocalMux I__1617 (
            .O(N__7189),
            .I(N__7186));
    Span4Mux_s3_h I__1616 (
            .O(N__7186),
            .I(N__7182));
    InMux I__1615 (
            .O(N__7185),
            .I(N__7179));
    Odrv4 I__1614 (
            .O(N__7182),
            .I(\uut.alu_out_m_0_2 ));
    LocalMux I__1613 (
            .O(N__7179),
            .I(\uut.alu_out_m_0_2 ));
    CascadeMux I__1612 (
            .O(N__7174),
            .I(\uut.out_1_0_iv_3_cascade_ ));
    CascadeMux I__1611 (
            .O(N__7171),
            .I(N__7168));
    InMux I__1610 (
            .O(N__7168),
            .I(N__7164));
    InMux I__1609 (
            .O(N__7167),
            .I(N__7160));
    LocalMux I__1608 (
            .O(N__7164),
            .I(N__7157));
    InMux I__1607 (
            .O(N__7163),
            .I(N__7154));
    LocalMux I__1606 (
            .O(N__7160),
            .I(N__7151));
    Span12Mux_s11_h I__1605 (
            .O(N__7157),
            .I(N__7148));
    LocalMux I__1604 (
            .O(N__7154),
            .I(\uut.AR_out_2 ));
    Odrv12 I__1603 (
            .O(N__7151),
            .I(\uut.AR_out_2 ));
    Odrv12 I__1602 (
            .O(N__7148),
            .I(\uut.AR_out_2 ));
    InMux I__1601 (
            .O(N__7141),
            .I(N__7136));
    InMux I__1600 (
            .O(N__7140),
            .I(N__7133));
    InMux I__1599 (
            .O(N__7139),
            .I(N__7129));
    LocalMux I__1598 (
            .O(N__7136),
            .I(N__7126));
    LocalMux I__1597 (
            .O(N__7133),
            .I(N__7123));
    InMux I__1596 (
            .O(N__7132),
            .I(N__7120));
    LocalMux I__1595 (
            .O(N__7129),
            .I(N__7117));
    Span4Mux_s2_h I__1594 (
            .O(N__7126),
            .I(N__7114));
    Span4Mux_v I__1593 (
            .O(N__7123),
            .I(N__7109));
    LocalMux I__1592 (
            .O(N__7120),
            .I(N__7109));
    Odrv4 I__1591 (
            .O(N__7117),
            .I(\uut.un11_MAR_LD ));
    Odrv4 I__1590 (
            .O(N__7114),
            .I(\uut.un11_MAR_LD ));
    Odrv4 I__1589 (
            .O(N__7109),
            .I(\uut.un11_MAR_LD ));
    InMux I__1588 (
            .O(N__7102),
            .I(N__7099));
    LocalMux I__1587 (
            .O(N__7099),
            .I(N__7096));
    Span4Mux_h I__1586 (
            .O(N__7096),
            .I(N__7093));
    Odrv4 I__1585 (
            .O(N__7093),
            .I(\uut.MAR_LD_1 ));
    InMux I__1584 (
            .O(N__7090),
            .I(N__7087));
    LocalMux I__1583 (
            .O(N__7087),
            .I(\uut.seq.counter.MAR_LD_0_0 ));
    CascadeMux I__1582 (
            .O(N__7084),
            .I(\uut.MAR_LD_1_cascade_ ));
    CascadeMux I__1581 (
            .O(N__7081),
            .I(N__7078));
    InMux I__1580 (
            .O(N__7078),
            .I(N__7075));
    LocalMux I__1579 (
            .O(N__7075),
            .I(\uut.N_16_0 ));
    InMux I__1578 (
            .O(N__7072),
            .I(N__7069));
    LocalMux I__1577 (
            .O(N__7069),
            .I(N__7066));
    Odrv4 I__1576 (
            .O(N__7066),
            .I(\uut.alu_out_m_1_3 ));
    CascadeMux I__1575 (
            .O(N__7063),
            .I(\uut.AR_BUF.g0Z0Z_5_cascade_ ));
    InMux I__1574 (
            .O(N__7060),
            .I(N__7056));
    CascadeMux I__1573 (
            .O(N__7059),
            .I(N__7053));
    LocalMux I__1572 (
            .O(N__7056),
            .I(N__7050));
    InMux I__1571 (
            .O(N__7053),
            .I(N__7046));
    Span4Mux_s2_h I__1570 (
            .O(N__7050),
            .I(N__7043));
    InMux I__1569 (
            .O(N__7049),
            .I(N__7040));
    LocalMux I__1568 (
            .O(N__7046),
            .I(\uut.seq.D_2_1 ));
    Odrv4 I__1567 (
            .O(N__7043),
            .I(\uut.seq.D_2_1 ));
    LocalMux I__1566 (
            .O(N__7040),
            .I(\uut.seq.D_2_1 ));
    InMux I__1565 (
            .O(N__7033),
            .I(N__7024));
    InMux I__1564 (
            .O(N__7032),
            .I(N__7021));
    CascadeMux I__1563 (
            .O(N__7031),
            .I(N__7016));
    CascadeMux I__1562 (
            .O(N__7030),
            .I(N__7013));
    InMux I__1561 (
            .O(N__7029),
            .I(N__7010));
    InMux I__1560 (
            .O(N__7028),
            .I(N__7007));
    InMux I__1559 (
            .O(N__7027),
            .I(N__7004));
    LocalMux I__1558 (
            .O(N__7024),
            .I(N__7001));
    LocalMux I__1557 (
            .O(N__7021),
            .I(N__6998));
    InMux I__1556 (
            .O(N__7020),
            .I(N__6995));
    InMux I__1555 (
            .O(N__7019),
            .I(N__6990));
    InMux I__1554 (
            .O(N__7016),
            .I(N__6990));
    InMux I__1553 (
            .O(N__7013),
            .I(N__6987));
    LocalMux I__1552 (
            .O(N__7010),
            .I(N__6982));
    LocalMux I__1551 (
            .O(N__7007),
            .I(N__6982));
    LocalMux I__1550 (
            .O(N__7004),
            .I(N__6979));
    Span4Mux_v I__1549 (
            .O(N__7001),
            .I(N__6976));
    Span12Mux_s4_h I__1548 (
            .O(N__6998),
            .I(N__6971));
    LocalMux I__1547 (
            .O(N__6995),
            .I(N__6971));
    LocalMux I__1546 (
            .O(N__6990),
            .I(N__6966));
    LocalMux I__1545 (
            .O(N__6987),
            .I(N__6966));
    Odrv4 I__1544 (
            .O(N__6982),
            .I(\uut.ir_out_i_2_6 ));
    Odrv12 I__1543 (
            .O(N__6979),
            .I(\uut.ir_out_i_2_6 ));
    Odrv4 I__1542 (
            .O(N__6976),
            .I(\uut.ir_out_i_2_6 ));
    Odrv12 I__1541 (
            .O(N__6971),
            .I(\uut.ir_out_i_2_6 ));
    Odrv4 I__1540 (
            .O(N__6966),
            .I(\uut.ir_out_i_2_6 ));
    CascadeMux I__1539 (
            .O(N__6955),
            .I(N__6952));
    InMux I__1538 (
            .O(N__6952),
            .I(N__6949));
    LocalMux I__1537 (
            .O(N__6949),
            .I(N__6946));
    Odrv4 I__1536 (
            .O(N__6946),
            .I(\uut.seq.D_2 ));
    InMux I__1535 (
            .O(N__6943),
            .I(N__6939));
    InMux I__1534 (
            .O(N__6942),
            .I(N__6936));
    LocalMux I__1533 (
            .O(N__6939),
            .I(N__6931));
    LocalMux I__1532 (
            .O(N__6936),
            .I(N__6928));
    InMux I__1531 (
            .O(N__6935),
            .I(N__6922));
    InMux I__1530 (
            .O(N__6934),
            .I(N__6919));
    Span4Mux_s3_h I__1529 (
            .O(N__6931),
            .I(N__6916));
    Span12Mux_s9_v I__1528 (
            .O(N__6928),
            .I(N__6913));
    InMux I__1527 (
            .O(N__6927),
            .I(N__6908));
    InMux I__1526 (
            .O(N__6926),
            .I(N__6908));
    InMux I__1525 (
            .O(N__6925),
            .I(N__6905));
    LocalMux I__1524 (
            .O(N__6922),
            .I(\uut.ir_out_i_2_5 ));
    LocalMux I__1523 (
            .O(N__6919),
            .I(\uut.ir_out_i_2_5 ));
    Odrv4 I__1522 (
            .O(N__6916),
            .I(\uut.ir_out_i_2_5 ));
    Odrv12 I__1521 (
            .O(N__6913),
            .I(\uut.ir_out_i_2_5 ));
    LocalMux I__1520 (
            .O(N__6908),
            .I(\uut.ir_out_i_2_5 ));
    LocalMux I__1519 (
            .O(N__6905),
            .I(\uut.ir_out_i_2_5 ));
    CascadeMux I__1518 (
            .O(N__6892),
            .I(\uut.B_LD_0_1_tz_cascade_ ));
    InMux I__1517 (
            .O(N__6889),
            .I(N__6886));
    LocalMux I__1516 (
            .O(N__6886),
            .I(N__6881));
    InMux I__1515 (
            .O(N__6885),
            .I(N__6878));
    CascadeMux I__1514 (
            .O(N__6884),
            .I(N__6875));
    Span4Mux_h I__1513 (
            .O(N__6881),
            .I(N__6869));
    LocalMux I__1512 (
            .O(N__6878),
            .I(N__6869));
    InMux I__1511 (
            .O(N__6875),
            .I(N__6866));
    InMux I__1510 (
            .O(N__6874),
            .I(N__6863));
    Span4Mux_h I__1509 (
            .O(N__6869),
            .I(N__6860));
    LocalMux I__1508 (
            .O(N__6866),
            .I(N__6857));
    LocalMux I__1507 (
            .O(N__6863),
            .I(N__6854));
    Odrv4 I__1506 (
            .O(N__6860),
            .I(\uut.mem.i2_mux_0 ));
    Odrv12 I__1505 (
            .O(N__6857),
            .I(\uut.mem.i2_mux_0 ));
    Odrv12 I__1504 (
            .O(N__6854),
            .I(\uut.mem.i2_mux_0 ));
    InMux I__1503 (
            .O(N__6847),
            .I(N__6844));
    LocalMux I__1502 (
            .O(N__6844),
            .I(N__6841));
    Odrv12 I__1501 (
            .O(N__6841),
            .I(\uut.out_1_0_iv_2_1 ));
    IoInMux I__1500 (
            .O(N__6838),
            .I(N__6835));
    LocalMux I__1499 (
            .O(N__6835),
            .I(N__6831));
    CascadeMux I__1498 (
            .O(N__6834),
            .I(N__6828));
    IoSpan4Mux I__1497 (
            .O(N__6831),
            .I(N__6825));
    InMux I__1496 (
            .O(N__6828),
            .I(N__6822));
    Odrv4 I__1495 (
            .O(N__6825),
            .I(LED3_c));
    LocalMux I__1494 (
            .O(N__6822),
            .I(LED3_c));
    InMux I__1493 (
            .O(N__6817),
            .I(N__6814));
    LocalMux I__1492 (
            .O(N__6814),
            .I(N__6811));
    Span4Mux_h I__1491 (
            .O(N__6811),
            .I(N__6808));
    Span4Mux_v I__1490 (
            .O(N__6808),
            .I(N__6805));
    Odrv4 I__1489 (
            .O(N__6805),
            .I(\uut.m10 ));
    CascadeMux I__1488 (
            .O(N__6802),
            .I(\uut.m10_cascade_ ));
    InMux I__1487 (
            .O(N__6799),
            .I(N__6795));
    InMux I__1486 (
            .O(N__6798),
            .I(N__6792));
    LocalMux I__1485 (
            .O(N__6795),
            .I(N__6789));
    LocalMux I__1484 (
            .O(N__6792),
            .I(N__6786));
    Span4Mux_s1_v I__1483 (
            .O(N__6789),
            .I(N__6783));
    Span4Mux_h I__1482 (
            .O(N__6786),
            .I(N__6780));
    Odrv4 I__1481 (
            .O(N__6783),
            .I(\uut.b_reg_out_0 ));
    Odrv4 I__1480 (
            .O(N__6780),
            .I(\uut.b_reg_out_0 ));
    InMux I__1479 (
            .O(N__6775),
            .I(N__6769));
    InMux I__1478 (
            .O(N__6774),
            .I(N__6763));
    InMux I__1477 (
            .O(N__6773),
            .I(N__6755));
    InMux I__1476 (
            .O(N__6772),
            .I(N__6755));
    LocalMux I__1475 (
            .O(N__6769),
            .I(N__6749));
    InMux I__1474 (
            .O(N__6768),
            .I(N__6746));
    InMux I__1473 (
            .O(N__6767),
            .I(N__6743));
    InMux I__1472 (
            .O(N__6766),
            .I(N__6740));
    LocalMux I__1471 (
            .O(N__6763),
            .I(N__6737));
    InMux I__1470 (
            .O(N__6762),
            .I(N__6732));
    InMux I__1469 (
            .O(N__6761),
            .I(N__6732));
    InMux I__1468 (
            .O(N__6760),
            .I(N__6729));
    LocalMux I__1467 (
            .O(N__6755),
            .I(N__6726));
    InMux I__1466 (
            .O(N__6754),
            .I(N__6723));
    InMux I__1465 (
            .O(N__6753),
            .I(N__6718));
    InMux I__1464 (
            .O(N__6752),
            .I(N__6718));
    Span4Mux_v I__1463 (
            .O(N__6749),
            .I(N__6713));
    LocalMux I__1462 (
            .O(N__6746),
            .I(N__6713));
    LocalMux I__1461 (
            .O(N__6743),
            .I(N__6706));
    LocalMux I__1460 (
            .O(N__6740),
            .I(N__6706));
    Span4Mux_v I__1459 (
            .O(N__6737),
            .I(N__6706));
    LocalMux I__1458 (
            .O(N__6732),
            .I(N__6703));
    LocalMux I__1457 (
            .O(N__6729),
            .I(N__6700));
    Span4Mux_s3_h I__1456 (
            .O(N__6726),
            .I(N__6693));
    LocalMux I__1455 (
            .O(N__6723),
            .I(N__6693));
    LocalMux I__1454 (
            .O(N__6718),
            .I(N__6693));
    Span4Mux_v I__1453 (
            .O(N__6713),
            .I(N__6690));
    Span4Mux_h I__1452 (
            .O(N__6706),
            .I(N__6685));
    Span4Mux_s2_h I__1451 (
            .O(N__6703),
            .I(N__6685));
    Span4Mux_h I__1450 (
            .O(N__6700),
            .I(N__6680));
    Span4Mux_v I__1449 (
            .O(N__6693),
            .I(N__6680));
    Odrv4 I__1448 (
            .O(N__6690),
            .I(\uut.T_1_fast_RNI28LI1_0 ));
    Odrv4 I__1447 (
            .O(N__6685),
            .I(\uut.T_1_fast_RNI28LI1_0 ));
    Odrv4 I__1446 (
            .O(N__6680),
            .I(\uut.T_1_fast_RNI28LI1_0 ));
    CascadeMux I__1445 (
            .O(N__6673),
            .I(N__6669));
    InMux I__1444 (
            .O(N__6672),
            .I(N__6665));
    InMux I__1443 (
            .O(N__6669),
            .I(N__6660));
    InMux I__1442 (
            .O(N__6668),
            .I(N__6660));
    LocalMux I__1441 (
            .O(N__6665),
            .I(N__6657));
    LocalMux I__1440 (
            .O(N__6660),
            .I(N__6654));
    Span4Mux_s2_h I__1439 (
            .O(N__6657),
            .I(N__6650));
    Span4Mux_s2_h I__1438 (
            .O(N__6654),
            .I(N__6647));
    InMux I__1437 (
            .O(N__6653),
            .I(N__6644));
    Odrv4 I__1436 (
            .O(N__6650),
            .I(\uut.b_reg_out_3 ));
    Odrv4 I__1435 (
            .O(N__6647),
            .I(\uut.b_reg_out_3 ));
    LocalMux I__1434 (
            .O(N__6644),
            .I(\uut.b_reg_out_3 ));
    InMux I__1433 (
            .O(N__6637),
            .I(N__6628));
    InMux I__1432 (
            .O(N__6636),
            .I(N__6628));
    InMux I__1431 (
            .O(N__6635),
            .I(N__6628));
    LocalMux I__1430 (
            .O(N__6628),
            .I(N__6625));
    Odrv4 I__1429 (
            .O(N__6625),
            .I(\uut.un1_A_cry_2_c_RNIBSP45 ));
    InMux I__1428 (
            .O(N__6622),
            .I(N__6611));
    InMux I__1427 (
            .O(N__6621),
            .I(N__6607));
    InMux I__1426 (
            .O(N__6620),
            .I(N__6604));
    InMux I__1425 (
            .O(N__6619),
            .I(N__6600));
    InMux I__1424 (
            .O(N__6618),
            .I(N__6597));
    InMux I__1423 (
            .O(N__6617),
            .I(N__6594));
    InMux I__1422 (
            .O(N__6616),
            .I(N__6591));
    InMux I__1421 (
            .O(N__6615),
            .I(N__6586));
    InMux I__1420 (
            .O(N__6614),
            .I(N__6586));
    LocalMux I__1419 (
            .O(N__6611),
            .I(N__6583));
    CascadeMux I__1418 (
            .O(N__6610),
            .I(N__6577));
    LocalMux I__1417 (
            .O(N__6607),
            .I(N__6572));
    LocalMux I__1416 (
            .O(N__6604),
            .I(N__6572));
    CascadeMux I__1415 (
            .O(N__6603),
            .I(N__6569));
    LocalMux I__1414 (
            .O(N__6600),
            .I(N__6566));
    LocalMux I__1413 (
            .O(N__6597),
            .I(N__6563));
    LocalMux I__1412 (
            .O(N__6594),
            .I(N__6560));
    LocalMux I__1411 (
            .O(N__6591),
            .I(N__6557));
    LocalMux I__1410 (
            .O(N__6586),
            .I(N__6554));
    Span4Mux_v I__1409 (
            .O(N__6583),
            .I(N__6551));
    InMux I__1408 (
            .O(N__6582),
            .I(N__6548));
    InMux I__1407 (
            .O(N__6581),
            .I(N__6543));
    InMux I__1406 (
            .O(N__6580),
            .I(N__6543));
    InMux I__1405 (
            .O(N__6577),
            .I(N__6540));
    Span4Mux_h I__1404 (
            .O(N__6572),
            .I(N__6537));
    InMux I__1403 (
            .O(N__6569),
            .I(N__6534));
    Span4Mux_h I__1402 (
            .O(N__6566),
            .I(N__6531));
    Span4Mux_v I__1401 (
            .O(N__6563),
            .I(N__6516));
    Span4Mux_v I__1400 (
            .O(N__6560),
            .I(N__6516));
    Span4Mux_h I__1399 (
            .O(N__6557),
            .I(N__6516));
    Span4Mux_v I__1398 (
            .O(N__6554),
            .I(N__6516));
    Span4Mux_s0_h I__1397 (
            .O(N__6551),
            .I(N__6516));
    LocalMux I__1396 (
            .O(N__6548),
            .I(N__6516));
    LocalMux I__1395 (
            .O(N__6543),
            .I(N__6516));
    LocalMux I__1394 (
            .O(N__6540),
            .I(\uut.un1_ALU_en_0 ));
    Odrv4 I__1393 (
            .O(N__6537),
            .I(\uut.un1_ALU_en_0 ));
    LocalMux I__1392 (
            .O(N__6534),
            .I(\uut.un1_ALU_en_0 ));
    Odrv4 I__1391 (
            .O(N__6531),
            .I(\uut.un1_ALU_en_0 ));
    Odrv4 I__1390 (
            .O(N__6516),
            .I(\uut.un1_ALU_en_0 ));
    CascadeMux I__1389 (
            .O(N__6505),
            .I(\uut.ALU_main.N_44_cascade_ ));
    InMux I__1388 (
            .O(N__6502),
            .I(N__6493));
    InMux I__1387 (
            .O(N__6501),
            .I(N__6489));
    InMux I__1386 (
            .O(N__6500),
            .I(N__6486));
    InMux I__1385 (
            .O(N__6499),
            .I(N__6479));
    InMux I__1384 (
            .O(N__6498),
            .I(N__6479));
    InMux I__1383 (
            .O(N__6497),
            .I(N__6479));
    CascadeMux I__1382 (
            .O(N__6496),
            .I(N__6476));
    LocalMux I__1381 (
            .O(N__6493),
            .I(N__6471));
    InMux I__1380 (
            .O(N__6492),
            .I(N__6468));
    LocalMux I__1379 (
            .O(N__6489),
            .I(N__6464));
    LocalMux I__1378 (
            .O(N__6486),
            .I(N__6460));
    LocalMux I__1377 (
            .O(N__6479),
            .I(N__6457));
    InMux I__1376 (
            .O(N__6476),
            .I(N__6453));
    InMux I__1375 (
            .O(N__6475),
            .I(N__6450));
    InMux I__1374 (
            .O(N__6474),
            .I(N__6447));
    Span4Mux_v I__1373 (
            .O(N__6471),
            .I(N__6442));
    LocalMux I__1372 (
            .O(N__6468),
            .I(N__6442));
    InMux I__1371 (
            .O(N__6467),
            .I(N__6439));
    Span4Mux_h I__1370 (
            .O(N__6464),
            .I(N__6436));
    InMux I__1369 (
            .O(N__6463),
            .I(N__6433));
    Span4Mux_v I__1368 (
            .O(N__6460),
            .I(N__6428));
    Span4Mux_v I__1367 (
            .O(N__6457),
            .I(N__6428));
    InMux I__1366 (
            .O(N__6456),
            .I(N__6425));
    LocalMux I__1365 (
            .O(N__6453),
            .I(\uut.T_1_fast_RNIVM0N3_0 ));
    LocalMux I__1364 (
            .O(N__6450),
            .I(\uut.T_1_fast_RNIVM0N3_0 ));
    LocalMux I__1363 (
            .O(N__6447),
            .I(\uut.T_1_fast_RNIVM0N3_0 ));
    Odrv4 I__1362 (
            .O(N__6442),
            .I(\uut.T_1_fast_RNIVM0N3_0 ));
    LocalMux I__1361 (
            .O(N__6439),
            .I(\uut.T_1_fast_RNIVM0N3_0 ));
    Odrv4 I__1360 (
            .O(N__6436),
            .I(\uut.T_1_fast_RNIVM0N3_0 ));
    LocalMux I__1359 (
            .O(N__6433),
            .I(\uut.T_1_fast_RNIVM0N3_0 ));
    Odrv4 I__1358 (
            .O(N__6428),
            .I(\uut.T_1_fast_RNIVM0N3_0 ));
    LocalMux I__1357 (
            .O(N__6425),
            .I(\uut.T_1_fast_RNIVM0N3_0 ));
    InMux I__1356 (
            .O(N__6406),
            .I(N__6403));
    LocalMux I__1355 (
            .O(N__6403),
            .I(N__6399));
    InMux I__1354 (
            .O(N__6402),
            .I(N__6396));
    Span4Mux_s1_h I__1353 (
            .O(N__6399),
            .I(N__6392));
    LocalMux I__1352 (
            .O(N__6396),
            .I(N__6389));
    InMux I__1351 (
            .O(N__6395),
            .I(N__6385));
    Span4Mux_h I__1350 (
            .O(N__6392),
            .I(N__6380));
    Span4Mux_h I__1349 (
            .O(N__6389),
            .I(N__6380));
    InMux I__1348 (
            .O(N__6388),
            .I(N__6377));
    LocalMux I__1347 (
            .O(N__6385),
            .I(N__6374));
    Odrv4 I__1346 (
            .O(N__6380),
            .I(\uut.acc_out_m_6 ));
    LocalMux I__1345 (
            .O(N__6377),
            .I(\uut.acc_out_m_6 ));
    Odrv12 I__1344 (
            .O(N__6374),
            .I(\uut.acc_out_m_6 ));
    InMux I__1343 (
            .O(N__6367),
            .I(N__6364));
    LocalMux I__1342 (
            .O(N__6364),
            .I(N__6360));
    InMux I__1341 (
            .O(N__6363),
            .I(N__6356));
    Span4Mux_v I__1340 (
            .O(N__6360),
            .I(N__6353));
    InMux I__1339 (
            .O(N__6359),
            .I(N__6350));
    LocalMux I__1338 (
            .O(N__6356),
            .I(N__6346));
    Span4Mux_h I__1337 (
            .O(N__6353),
            .I(N__6341));
    LocalMux I__1336 (
            .O(N__6350),
            .I(N__6341));
    InMux I__1335 (
            .O(N__6349),
            .I(N__6338));
    Odrv4 I__1334 (
            .O(N__6346),
            .I(\uut.alu_out_m_6 ));
    Odrv4 I__1333 (
            .O(N__6341),
            .I(\uut.alu_out_m_6 ));
    LocalMux I__1332 (
            .O(N__6338),
            .I(\uut.alu_out_m_6 ));
    CascadeMux I__1331 (
            .O(N__6331),
            .I(N__6327));
    CascadeMux I__1330 (
            .O(N__6330),
            .I(N__6324));
    InMux I__1329 (
            .O(N__6327),
            .I(N__6321));
    InMux I__1328 (
            .O(N__6324),
            .I(N__6317));
    LocalMux I__1327 (
            .O(N__6321),
            .I(N__6313));
    CascadeMux I__1326 (
            .O(N__6320),
            .I(N__6310));
    LocalMux I__1325 (
            .O(N__6317),
            .I(N__6307));
    CascadeMux I__1324 (
            .O(N__6316),
            .I(N__6304));
    Span4Mux_v I__1323 (
            .O(N__6313),
            .I(N__6301));
    InMux I__1322 (
            .O(N__6310),
            .I(N__6298));
    Span4Mux_v I__1321 (
            .O(N__6307),
            .I(N__6295));
    InMux I__1320 (
            .O(N__6304),
            .I(N__6292));
    Span4Mux_h I__1319 (
            .O(N__6301),
            .I(N__6289));
    LocalMux I__1318 (
            .O(N__6298),
            .I(N__6286));
    Sp12to4 I__1317 (
            .O(N__6295),
            .I(N__6281));
    LocalMux I__1316 (
            .O(N__6292),
            .I(N__6281));
    Odrv4 I__1315 (
            .O(N__6289),
            .I(\uut.mem.N_29_mux ));
    Odrv4 I__1314 (
            .O(N__6286),
            .I(\uut.mem.N_29_mux ));
    Odrv12 I__1313 (
            .O(N__6281),
            .I(\uut.mem.N_29_mux ));
    CascadeMux I__1312 (
            .O(N__6274),
            .I(N__6269));
    InMux I__1311 (
            .O(N__6273),
            .I(N__6266));
    InMux I__1310 (
            .O(N__6272),
            .I(N__6262));
    InMux I__1309 (
            .O(N__6269),
            .I(N__6259));
    LocalMux I__1308 (
            .O(N__6266),
            .I(N__6256));
    InMux I__1307 (
            .O(N__6265),
            .I(N__6253));
    LocalMux I__1306 (
            .O(N__6262),
            .I(N__6250));
    LocalMux I__1305 (
            .O(N__6259),
            .I(N__6247));
    Span4Mux_h I__1304 (
            .O(N__6256),
            .I(N__6244));
    LocalMux I__1303 (
            .O(N__6253),
            .I(N__6239));
    Span12Mux_v I__1302 (
            .O(N__6250),
            .I(N__6239));
    Span4Mux_v I__1301 (
            .O(N__6247),
            .I(N__6236));
    Odrv4 I__1300 (
            .O(N__6244),
            .I(\uut.acc_out_6 ));
    Odrv12 I__1299 (
            .O(N__6239),
            .I(\uut.acc_out_6 ));
    Odrv4 I__1298 (
            .O(N__6236),
            .I(\uut.acc_out_6 ));
    CascadeMux I__1297 (
            .O(N__6229),
            .I(N__6225));
    InMux I__1296 (
            .O(N__6228),
            .I(N__6222));
    InMux I__1295 (
            .O(N__6225),
            .I(N__6219));
    LocalMux I__1294 (
            .O(N__6222),
            .I(N__6216));
    LocalMux I__1293 (
            .O(N__6219),
            .I(N__6210));
    Span4Mux_s1_h I__1292 (
            .O(N__6216),
            .I(N__6210));
    InMux I__1291 (
            .O(N__6215),
            .I(N__6207));
    Span4Mux_h I__1290 (
            .O(N__6210),
            .I(N__6204));
    LocalMux I__1289 (
            .O(N__6207),
            .I(\uut.acc_out_m_7 ));
    Odrv4 I__1288 (
            .O(N__6204),
            .I(\uut.acc_out_m_7 ));
    InMux I__1287 (
            .O(N__6199),
            .I(N__6196));
    LocalMux I__1286 (
            .O(N__6196),
            .I(N__6191));
    InMux I__1285 (
            .O(N__6195),
            .I(N__6188));
    InMux I__1284 (
            .O(N__6194),
            .I(N__6185));
    Odrv12 I__1283 (
            .O(N__6191),
            .I(\uut.alu_out_m_7 ));
    LocalMux I__1282 (
            .O(N__6188),
            .I(\uut.alu_out_m_7 ));
    LocalMux I__1281 (
            .O(N__6185),
            .I(\uut.alu_out_m_7 ));
    InMux I__1280 (
            .O(N__6178),
            .I(N__6174));
    InMux I__1279 (
            .O(N__6177),
            .I(N__6171));
    LocalMux I__1278 (
            .O(N__6174),
            .I(N__6165));
    LocalMux I__1277 (
            .O(N__6171),
            .I(N__6165));
    InMux I__1276 (
            .O(N__6170),
            .I(N__6162));
    Span4Mux_s3_v I__1275 (
            .O(N__6165),
            .I(N__6159));
    LocalMux I__1274 (
            .O(N__6162),
            .I(N__6156));
    Span4Mux_h I__1273 (
            .O(N__6159),
            .I(N__6153));
    Span4Mux_h I__1272 (
            .O(N__6156),
            .I(N__6150));
    Odrv4 I__1271 (
            .O(N__6153),
            .I(\uut.acc_out_7 ));
    Odrv4 I__1270 (
            .O(N__6150),
            .I(\uut.acc_out_7 ));
    InMux I__1269 (
            .O(N__6145),
            .I(N__6142));
    LocalMux I__1268 (
            .O(N__6142),
            .I(N__6138));
    InMux I__1267 (
            .O(N__6141),
            .I(N__6135));
    Span4Mux_v I__1266 (
            .O(N__6138),
            .I(N__6132));
    LocalMux I__1265 (
            .O(N__6135),
            .I(N__6129));
    Span4Mux_h I__1264 (
            .O(N__6132),
            .I(N__6123));
    Span4Mux_v I__1263 (
            .O(N__6129),
            .I(N__6123));
    InMux I__1262 (
            .O(N__6128),
            .I(N__6120));
    Odrv4 I__1261 (
            .O(N__6123),
            .I(\uut.alu_out_m_5 ));
    LocalMux I__1260 (
            .O(N__6120),
            .I(\uut.alu_out_m_5 ));
    InMux I__1259 (
            .O(N__6115),
            .I(N__6111));
    InMux I__1258 (
            .O(N__6114),
            .I(N__6108));
    LocalMux I__1257 (
            .O(N__6111),
            .I(N__6105));
    LocalMux I__1256 (
            .O(N__6108),
            .I(N__6102));
    Span12Mux_s6_h I__1255 (
            .O(N__6105),
            .I(N__6097));
    Span4Mux_v I__1254 (
            .O(N__6102),
            .I(N__6094));
    InMux I__1253 (
            .O(N__6101),
            .I(N__6091));
    InMux I__1252 (
            .O(N__6100),
            .I(N__6088));
    Odrv12 I__1251 (
            .O(N__6097),
            .I(\uut.acc_out_m_5 ));
    Odrv4 I__1250 (
            .O(N__6094),
            .I(\uut.acc_out_m_5 ));
    LocalMux I__1249 (
            .O(N__6091),
            .I(\uut.acc_out_m_5 ));
    LocalMux I__1248 (
            .O(N__6088),
            .I(\uut.acc_out_m_5 ));
    CascadeMux I__1247 (
            .O(N__6079),
            .I(N__6075));
    InMux I__1246 (
            .O(N__6078),
            .I(N__6071));
    InMux I__1245 (
            .O(N__6075),
            .I(N__6067));
    InMux I__1244 (
            .O(N__6074),
            .I(N__6064));
    LocalMux I__1243 (
            .O(N__6071),
            .I(N__6061));
    CascadeMux I__1242 (
            .O(N__6070),
            .I(N__6058));
    LocalMux I__1241 (
            .O(N__6067),
            .I(N__6053));
    LocalMux I__1240 (
            .O(N__6064),
            .I(N__6053));
    Span4Mux_h I__1239 (
            .O(N__6061),
            .I(N__6050));
    InMux I__1238 (
            .O(N__6058),
            .I(N__6047));
    Span4Mux_h I__1237 (
            .O(N__6053),
            .I(N__6044));
    Sp12to4 I__1236 (
            .O(N__6050),
            .I(N__6039));
    LocalMux I__1235 (
            .O(N__6047),
            .I(N__6039));
    Span4Mux_h I__1234 (
            .O(N__6044),
            .I(N__6036));
    Odrv12 I__1233 (
            .O(N__6039),
            .I(\uut.mem.m20 ));
    Odrv4 I__1232 (
            .O(N__6036),
            .I(\uut.mem.m20 ));
    CascadeMux I__1231 (
            .O(N__6031),
            .I(N__6025));
    InMux I__1230 (
            .O(N__6030),
            .I(N__6022));
    InMux I__1229 (
            .O(N__6029),
            .I(N__6019));
    CascadeMux I__1228 (
            .O(N__6028),
            .I(N__6016));
    InMux I__1227 (
            .O(N__6025),
            .I(N__6013));
    LocalMux I__1226 (
            .O(N__6022),
            .I(N__6010));
    LocalMux I__1225 (
            .O(N__6019),
            .I(N__6007));
    InMux I__1224 (
            .O(N__6016),
            .I(N__6004));
    LocalMux I__1223 (
            .O(N__6013),
            .I(N__6001));
    Span4Mux_v I__1222 (
            .O(N__6010),
            .I(N__5994));
    Span4Mux_h I__1221 (
            .O(N__6007),
            .I(N__5994));
    LocalMux I__1220 (
            .O(N__6004),
            .I(N__5994));
    Span4Mux_h I__1219 (
            .O(N__6001),
            .I(N__5991));
    Span4Mux_h I__1218 (
            .O(N__5994),
            .I(N__5988));
    Odrv4 I__1217 (
            .O(N__5991),
            .I(\uut.acc_out_5 ));
    Odrv4 I__1216 (
            .O(N__5988),
            .I(\uut.acc_out_5 ));
    CascadeMux I__1215 (
            .O(N__5983),
            .I(N__5980));
    InMux I__1214 (
            .O(N__5980),
            .I(N__5976));
    InMux I__1213 (
            .O(N__5979),
            .I(N__5973));
    LocalMux I__1212 (
            .O(N__5976),
            .I(N__5970));
    LocalMux I__1211 (
            .O(N__5973),
            .I(N__5967));
    Span4Mux_v I__1210 (
            .O(N__5970),
            .I(N__5961));
    Span4Mux_v I__1209 (
            .O(N__5967),
            .I(N__5961));
    InMux I__1208 (
            .O(N__5966),
            .I(N__5958));
    Odrv4 I__1207 (
            .O(N__5961),
            .I(\uut.q_RNIDGA71 ));
    LocalMux I__1206 (
            .O(N__5958),
            .I(\uut.q_RNIDGA71 ));
    CascadeMux I__1205 (
            .O(N__5953),
            .I(N__5950));
    InMux I__1204 (
            .O(N__5950),
            .I(N__5943));
    InMux I__1203 (
            .O(N__5949),
            .I(N__5940));
    InMux I__1202 (
            .O(N__5948),
            .I(N__5933));
    InMux I__1201 (
            .O(N__5947),
            .I(N__5933));
    InMux I__1200 (
            .O(N__5946),
            .I(N__5933));
    LocalMux I__1199 (
            .O(N__5943),
            .I(N__5930));
    LocalMux I__1198 (
            .O(N__5940),
            .I(N__5925));
    LocalMux I__1197 (
            .O(N__5933),
            .I(N__5925));
    Span4Mux_v I__1196 (
            .O(N__5930),
            .I(N__5920));
    Span4Mux_v I__1195 (
            .O(N__5925),
            .I(N__5920));
    Odrv4 I__1194 (
            .O(N__5920),
            .I(\uut.mem.i2_mux ));
    InMux I__1193 (
            .O(N__5917),
            .I(N__5914));
    LocalMux I__1192 (
            .O(N__5914),
            .I(N__5910));
    InMux I__1191 (
            .O(N__5913),
            .I(N__5907));
    Span4Mux_v I__1190 (
            .O(N__5910),
            .I(N__5902));
    LocalMux I__1189 (
            .O(N__5907),
            .I(N__5899));
    InMux I__1188 (
            .O(N__5906),
            .I(N__5896));
    InMux I__1187 (
            .O(N__5905),
            .I(N__5893));
    Odrv4 I__1186 (
            .O(N__5902),
            .I(\uut.alu_out_m_4 ));
    Odrv4 I__1185 (
            .O(N__5899),
            .I(\uut.alu_out_m_4 ));
    LocalMux I__1184 (
            .O(N__5896),
            .I(\uut.alu_out_m_4 ));
    LocalMux I__1183 (
            .O(N__5893),
            .I(\uut.alu_out_m_4 ));
    CascadeMux I__1182 (
            .O(N__5884),
            .I(N__5880));
    CascadeMux I__1181 (
            .O(N__5883),
            .I(N__5874));
    InMux I__1180 (
            .O(N__5880),
            .I(N__5871));
    InMux I__1179 (
            .O(N__5879),
            .I(N__5864));
    InMux I__1178 (
            .O(N__5878),
            .I(N__5864));
    InMux I__1177 (
            .O(N__5877),
            .I(N__5864));
    InMux I__1176 (
            .O(N__5874),
            .I(N__5861));
    LocalMux I__1175 (
            .O(N__5871),
            .I(N__5856));
    LocalMux I__1174 (
            .O(N__5864),
            .I(N__5856));
    LocalMux I__1173 (
            .O(N__5861),
            .I(N__5853));
    Span4Mux_h I__1172 (
            .O(N__5856),
            .I(N__5848));
    Span4Mux_h I__1171 (
            .O(N__5853),
            .I(N__5848));
    Odrv4 I__1170 (
            .O(N__5848),
            .I(\uut.acc_out_4 ));
    CEMux I__1169 (
            .O(N__5845),
            .I(N__5842));
    LocalMux I__1168 (
            .O(N__5842),
            .I(N__5838));
    CEMux I__1167 (
            .O(N__5841),
            .I(N__5834));
    Span4Mux_h I__1166 (
            .O(N__5838),
            .I(N__5830));
    CEMux I__1165 (
            .O(N__5837),
            .I(N__5827));
    LocalMux I__1164 (
            .O(N__5834),
            .I(N__5824));
    CEMux I__1163 (
            .O(N__5833),
            .I(N__5821));
    Span4Mux_v I__1162 (
            .O(N__5830),
            .I(N__5816));
    LocalMux I__1161 (
            .O(N__5827),
            .I(N__5816));
    Span4Mux_v I__1160 (
            .O(N__5824),
            .I(N__5813));
    LocalMux I__1159 (
            .O(N__5821),
            .I(N__5810));
    Span4Mux_s3_h I__1158 (
            .O(N__5816),
            .I(N__5807));
    Span4Mux_h I__1157 (
            .O(N__5813),
            .I(N__5802));
    Span4Mux_v I__1156 (
            .O(N__5810),
            .I(N__5802));
    Odrv4 I__1155 (
            .O(N__5807),
            .I(\uut.ACC_LD_0_i ));
    Odrv4 I__1154 (
            .O(N__5802),
            .I(\uut.ACC_LD_0_i ));
    InMux I__1153 (
            .O(N__5797),
            .I(N__5794));
    LocalMux I__1152 (
            .O(N__5794),
            .I(N__5789));
    InMux I__1151 (
            .O(N__5793),
            .I(N__5786));
    CascadeMux I__1150 (
            .O(N__5792),
            .I(N__5783));
    Span4Mux_h I__1149 (
            .O(N__5789),
            .I(N__5780));
    LocalMux I__1148 (
            .O(N__5786),
            .I(N__5777));
    InMux I__1147 (
            .O(N__5783),
            .I(N__5774));
    Odrv4 I__1146 (
            .O(N__5780),
            .I(\uut.program_counter_2 ));
    Odrv12 I__1145 (
            .O(N__5777),
            .I(\uut.program_counter_2 ));
    LocalMux I__1144 (
            .O(N__5774),
            .I(\uut.program_counter_2 ));
    CascadeMux I__1143 (
            .O(N__5767),
            .I(N__5764));
    InMux I__1142 (
            .O(N__5764),
            .I(N__5760));
    CascadeMux I__1141 (
            .O(N__5763),
            .I(N__5757));
    LocalMux I__1140 (
            .O(N__5760),
            .I(N__5754));
    InMux I__1139 (
            .O(N__5757),
            .I(N__5751));
    Span4Mux_v I__1138 (
            .O(N__5754),
            .I(N__5745));
    LocalMux I__1137 (
            .O(N__5751),
            .I(N__5742));
    InMux I__1136 (
            .O(N__5750),
            .I(N__5739));
    CascadeMux I__1135 (
            .O(N__5749),
            .I(N__5736));
    CascadeMux I__1134 (
            .O(N__5748),
            .I(N__5733));
    Span4Mux_h I__1133 (
            .O(N__5745),
            .I(N__5730));
    Span4Mux_s2_h I__1132 (
            .O(N__5742),
            .I(N__5725));
    LocalMux I__1131 (
            .O(N__5739),
            .I(N__5725));
    InMux I__1130 (
            .O(N__5736),
            .I(N__5720));
    InMux I__1129 (
            .O(N__5733),
            .I(N__5720));
    Odrv4 I__1128 (
            .O(N__5730),
            .I(\uut.program_counter_1 ));
    Odrv4 I__1127 (
            .O(N__5725),
            .I(\uut.program_counter_1 ));
    LocalMux I__1126 (
            .O(N__5720),
            .I(\uut.program_counter_1 ));
    InMux I__1125 (
            .O(N__5713),
            .I(N__5710));
    LocalMux I__1124 (
            .O(N__5710),
            .I(N__5706));
    InMux I__1123 (
            .O(N__5709),
            .I(N__5703));
    Span4Mux_s3_h I__1122 (
            .O(N__5706),
            .I(N__5697));
    LocalMux I__1121 (
            .O(N__5703),
            .I(N__5694));
    InMux I__1120 (
            .O(N__5702),
            .I(N__5687));
    InMux I__1119 (
            .O(N__5701),
            .I(N__5687));
    InMux I__1118 (
            .O(N__5700),
            .I(N__5687));
    Odrv4 I__1117 (
            .O(N__5697),
            .I(\uut.program_counter_0 ));
    Odrv12 I__1116 (
            .O(N__5694),
            .I(\uut.program_counter_0 ));
    LocalMux I__1115 (
            .O(N__5687),
            .I(\uut.program_counter_0 ));
    InMux I__1114 (
            .O(N__5680),
            .I(N__5677));
    LocalMux I__1113 (
            .O(N__5677),
            .I(\uut.pc.program_counter_RNO_1Z0Z_2 ));
    CascadeMux I__1112 (
            .O(N__5674),
            .I(\uut.N_44_0_cascade_ ));
    InMux I__1111 (
            .O(N__5671),
            .I(N__5668));
    LocalMux I__1110 (
            .O(N__5668),
            .I(N__5665));
    Odrv4 I__1109 (
            .O(N__5665),
            .I(\uut.pc.g0_rn_1 ));
    CascadeMux I__1108 (
            .O(N__5662),
            .I(\uut.pc.alu_out_m_0_3_cascade_ ));
    ClkMux I__1107 (
            .O(N__5659),
            .I(N__5548));
    ClkMux I__1106 (
            .O(N__5658),
            .I(N__5548));
    ClkMux I__1105 (
            .O(N__5657),
            .I(N__5548));
    ClkMux I__1104 (
            .O(N__5656),
            .I(N__5548));
    ClkMux I__1103 (
            .O(N__5655),
            .I(N__5548));
    ClkMux I__1102 (
            .O(N__5654),
            .I(N__5548));
    ClkMux I__1101 (
            .O(N__5653),
            .I(N__5548));
    ClkMux I__1100 (
            .O(N__5652),
            .I(N__5548));
    ClkMux I__1099 (
            .O(N__5651),
            .I(N__5548));
    ClkMux I__1098 (
            .O(N__5650),
            .I(N__5548));
    ClkMux I__1097 (
            .O(N__5649),
            .I(N__5548));
    ClkMux I__1096 (
            .O(N__5648),
            .I(N__5548));
    ClkMux I__1095 (
            .O(N__5647),
            .I(N__5548));
    ClkMux I__1094 (
            .O(N__5646),
            .I(N__5548));
    ClkMux I__1093 (
            .O(N__5645),
            .I(N__5548));
    ClkMux I__1092 (
            .O(N__5644),
            .I(N__5548));
    ClkMux I__1091 (
            .O(N__5643),
            .I(N__5548));
    ClkMux I__1090 (
            .O(N__5642),
            .I(N__5548));
    ClkMux I__1089 (
            .O(N__5641),
            .I(N__5548));
    ClkMux I__1088 (
            .O(N__5640),
            .I(N__5548));
    ClkMux I__1087 (
            .O(N__5639),
            .I(N__5548));
    ClkMux I__1086 (
            .O(N__5638),
            .I(N__5548));
    ClkMux I__1085 (
            .O(N__5637),
            .I(N__5548));
    ClkMux I__1084 (
            .O(N__5636),
            .I(N__5548));
    ClkMux I__1083 (
            .O(N__5635),
            .I(N__5548));
    ClkMux I__1082 (
            .O(N__5634),
            .I(N__5548));
    ClkMux I__1081 (
            .O(N__5633),
            .I(N__5548));
    ClkMux I__1080 (
            .O(N__5632),
            .I(N__5548));
    ClkMux I__1079 (
            .O(N__5631),
            .I(N__5548));
    ClkMux I__1078 (
            .O(N__5630),
            .I(N__5548));
    ClkMux I__1077 (
            .O(N__5629),
            .I(N__5548));
    ClkMux I__1076 (
            .O(N__5628),
            .I(N__5548));
    ClkMux I__1075 (
            .O(N__5627),
            .I(N__5548));
    ClkMux I__1074 (
            .O(N__5626),
            .I(N__5548));
    ClkMux I__1073 (
            .O(N__5625),
            .I(N__5548));
    ClkMux I__1072 (
            .O(N__5624),
            .I(N__5548));
    ClkMux I__1071 (
            .O(N__5623),
            .I(N__5548));
    GlobalMux I__1070 (
            .O(N__5548),
            .I(N__5545));
    gio2CtrlBuf I__1069 (
            .O(N__5545),
            .I(\uut.buf_clk_1_g ));
    CascadeMux I__1068 (
            .O(N__5542),
            .I(N__5539));
    InMux I__1067 (
            .O(N__5539),
            .I(N__5536));
    LocalMux I__1066 (
            .O(N__5536),
            .I(N__5533));
    Odrv4 I__1065 (
            .O(N__5533),
            .I(\uut.ALU_main.N_44_1 ));
    InMux I__1064 (
            .O(N__5530),
            .I(N__5527));
    LocalMux I__1063 (
            .O(N__5527),
            .I(\uut.pc.g1 ));
    CascadeMux I__1062 (
            .O(N__5524),
            .I(\uut.pc.un1_inc_0_0_cascade_ ));
    InMux I__1061 (
            .O(N__5521),
            .I(N__5517));
    InMux I__1060 (
            .O(N__5520),
            .I(N__5513));
    LocalMux I__1059 (
            .O(N__5517),
            .I(N__5510));
    InMux I__1058 (
            .O(N__5516),
            .I(N__5507));
    LocalMux I__1057 (
            .O(N__5513),
            .I(N__5502));
    Span4Mux_s3_h I__1056 (
            .O(N__5510),
            .I(N__5502));
    LocalMux I__1055 (
            .O(N__5507),
            .I(N__5499));
    Odrv4 I__1054 (
            .O(N__5502),
            .I(\uut.un17_IR_OE ));
    Odrv12 I__1053 (
            .O(N__5499),
            .I(\uut.un17_IR_OE ));
    InMux I__1052 (
            .O(N__5494),
            .I(N__5491));
    LocalMux I__1051 (
            .O(N__5491),
            .I(\uut.PC_LD_0_0 ));
    CascadeMux I__1050 (
            .O(N__5488),
            .I(\uut.PC_LD_0_0_cascade_ ));
    InMux I__1049 (
            .O(N__5485),
            .I(N__5481));
    CascadeMux I__1048 (
            .O(N__5484),
            .I(N__5478));
    LocalMux I__1047 (
            .O(N__5481),
            .I(N__5475));
    InMux I__1046 (
            .O(N__5478),
            .I(N__5472));
    Span4Mux_v I__1045 (
            .O(N__5475),
            .I(N__5467));
    LocalMux I__1044 (
            .O(N__5472),
            .I(N__5467));
    Odrv4 I__1043 (
            .O(N__5467),
            .I(\uut.pc.un1_inc_0 ));
    CascadeMux I__1042 (
            .O(N__5464),
            .I(\uut.pc.un1_inc_0_cascade_ ));
    InMux I__1041 (
            .O(N__5461),
            .I(N__5458));
    LocalMux I__1040 (
            .O(N__5458),
            .I(N__5455));
    Odrv12 I__1039 (
            .O(N__5455),
            .I(\uut.pc.program_counter_4_1_2 ));
    CascadeMux I__1038 (
            .O(N__5452),
            .I(N__5448));
    CascadeMux I__1037 (
            .O(N__5451),
            .I(N__5445));
    InMux I__1036 (
            .O(N__5448),
            .I(N__5442));
    InMux I__1035 (
            .O(N__5445),
            .I(N__5439));
    LocalMux I__1034 (
            .O(N__5442),
            .I(N__5436));
    LocalMux I__1033 (
            .O(N__5439),
            .I(N__5433));
    Span12Mux_s10_v I__1032 (
            .O(N__5436),
            .I(N__5430));
    Span4Mux_h I__1031 (
            .O(N__5433),
            .I(N__5427));
    Odrv12 I__1030 (
            .O(N__5430),
            .I(\uut.m13 ));
    Odrv4 I__1029 (
            .O(N__5427),
            .I(\uut.m13 ));
    InMux I__1028 (
            .O(N__5422),
            .I(N__5410));
    InMux I__1027 (
            .O(N__5421),
            .I(N__5407));
    InMux I__1026 (
            .O(N__5420),
            .I(N__5402));
    InMux I__1025 (
            .O(N__5419),
            .I(N__5402));
    InMux I__1024 (
            .O(N__5418),
            .I(N__5395));
    InMux I__1023 (
            .O(N__5417),
            .I(N__5395));
    InMux I__1022 (
            .O(N__5416),
            .I(N__5395));
    InMux I__1021 (
            .O(N__5415),
            .I(N__5388));
    InMux I__1020 (
            .O(N__5414),
            .I(N__5388));
    InMux I__1019 (
            .O(N__5413),
            .I(N__5388));
    LocalMux I__1018 (
            .O(N__5410),
            .I(\uut.q_0_fast_0 ));
    LocalMux I__1017 (
            .O(N__5407),
            .I(\uut.q_0_fast_0 ));
    LocalMux I__1016 (
            .O(N__5402),
            .I(\uut.q_0_fast_0 ));
    LocalMux I__1015 (
            .O(N__5395),
            .I(\uut.q_0_fast_0 ));
    LocalMux I__1014 (
            .O(N__5388),
            .I(\uut.q_0_fast_0 ));
    CascadeMux I__1013 (
            .O(N__5377),
            .I(N__5373));
    InMux I__1012 (
            .O(N__5376),
            .I(N__5370));
    InMux I__1011 (
            .O(N__5373),
            .I(N__5367));
    LocalMux I__1010 (
            .O(N__5370),
            .I(\uut.seq.counter.T_fastZ0Z_2 ));
    LocalMux I__1009 (
            .O(N__5367),
            .I(\uut.seq.counter.T_fastZ0Z_2 ));
    CascadeMux I__1008 (
            .O(N__5362),
            .I(\uut.seq.counter.T_fast_RNIH09PZ0Z_2_cascade_ ));
    InMux I__1007 (
            .O(N__5359),
            .I(N__5353));
    CascadeMux I__1006 (
            .O(N__5358),
            .I(N__5350));
    InMux I__1005 (
            .O(N__5357),
            .I(N__5346));
    CascadeMux I__1004 (
            .O(N__5356),
            .I(N__5343));
    LocalMux I__1003 (
            .O(N__5353),
            .I(N__5336));
    InMux I__1002 (
            .O(N__5350),
            .I(N__5331));
    InMux I__1001 (
            .O(N__5349),
            .I(N__5331));
    LocalMux I__1000 (
            .O(N__5346),
            .I(N__5328));
    InMux I__999 (
            .O(N__5343),
            .I(N__5325));
    InMux I__998 (
            .O(N__5342),
            .I(N__5322));
    InMux I__997 (
            .O(N__5341),
            .I(N__5315));
    InMux I__996 (
            .O(N__5340),
            .I(N__5315));
    InMux I__995 (
            .O(N__5339),
            .I(N__5315));
    Odrv4 I__994 (
            .O(N__5336),
            .I(\uut.ir_out_4_rep1 ));
    LocalMux I__993 (
            .O(N__5331),
            .I(\uut.ir_out_4_rep1 ));
    Odrv12 I__992 (
            .O(N__5328),
            .I(\uut.ir_out_4_rep1 ));
    LocalMux I__991 (
            .O(N__5325),
            .I(\uut.ir_out_4_rep1 ));
    LocalMux I__990 (
            .O(N__5322),
            .I(\uut.ir_out_4_rep1 ));
    LocalMux I__989 (
            .O(N__5315),
            .I(\uut.ir_out_4_rep1 ));
    InMux I__988 (
            .O(N__5302),
            .I(N__5294));
    InMux I__987 (
            .O(N__5301),
            .I(N__5289));
    InMux I__986 (
            .O(N__5300),
            .I(N__5289));
    InMux I__985 (
            .O(N__5299),
            .I(N__5284));
    InMux I__984 (
            .O(N__5298),
            .I(N__5284));
    InMux I__983 (
            .O(N__5297),
            .I(N__5280));
    LocalMux I__982 (
            .O(N__5294),
            .I(N__5277));
    LocalMux I__981 (
            .O(N__5289),
            .I(N__5272));
    LocalMux I__980 (
            .O(N__5284),
            .I(N__5272));
    InMux I__979 (
            .O(N__5283),
            .I(N__5269));
    LocalMux I__978 (
            .O(N__5280),
            .I(N__5266));
    Span4Mux_h I__977 (
            .O(N__5277),
            .I(N__5261));
    Span4Mux_v I__976 (
            .O(N__5272),
            .I(N__5261));
    LocalMux I__975 (
            .O(N__5269),
            .I(N__5258));
    Span4Mux_v I__974 (
            .O(N__5266),
            .I(N__5255));
    Span4Mux_v I__973 (
            .O(N__5261),
            .I(N__5250));
    Span4Mux_s1_v I__972 (
            .O(N__5258),
            .I(N__5250));
    Odrv4 I__971 (
            .O(N__5255),
            .I(\uut.ir_out_0 ));
    Odrv4 I__970 (
            .O(N__5250),
            .I(\uut.ir_out_0 ));
    CascadeMux I__969 (
            .O(N__5245),
            .I(N__5238));
    InMux I__968 (
            .O(N__5244),
            .I(N__5234));
    InMux I__967 (
            .O(N__5243),
            .I(N__5231));
    InMux I__966 (
            .O(N__5242),
            .I(N__5226));
    InMux I__965 (
            .O(N__5241),
            .I(N__5226));
    InMux I__964 (
            .O(N__5238),
            .I(N__5221));
    InMux I__963 (
            .O(N__5237),
            .I(N__5221));
    LocalMux I__962 (
            .O(N__5234),
            .I(N__5214));
    LocalMux I__961 (
            .O(N__5231),
            .I(N__5214));
    LocalMux I__960 (
            .O(N__5226),
            .I(N__5214));
    LocalMux I__959 (
            .O(N__5221),
            .I(\uut.acc_out_0 ));
    Odrv12 I__958 (
            .O(N__5214),
            .I(\uut.acc_out_0 ));
    CascadeMux I__957 (
            .O(N__5209),
            .I(\uut.OUT_LD_cascade_ ));
    InMux I__956 (
            .O(N__5206),
            .I(N__5203));
    LocalMux I__955 (
            .O(N__5203),
            .I(N__5200));
    Span4Mux_v I__954 (
            .O(N__5200),
            .I(N__5197));
    Odrv4 I__953 (
            .O(N__5197),
            .I(\uut.pc.G_26_i_a4_1 ));
    CascadeMux I__952 (
            .O(N__5194),
            .I(N__5189));
    CascadeMux I__951 (
            .O(N__5193),
            .I(N__5186));
    CascadeMux I__950 (
            .O(N__5192),
            .I(N__5183));
    InMux I__949 (
            .O(N__5189),
            .I(N__5178));
    InMux I__948 (
            .O(N__5186),
            .I(N__5175));
    InMux I__947 (
            .O(N__5183),
            .I(N__5172));
    InMux I__946 (
            .O(N__5182),
            .I(N__5168));
    InMux I__945 (
            .O(N__5181),
            .I(N__5165));
    LocalMux I__944 (
            .O(N__5178),
            .I(N__5160));
    LocalMux I__943 (
            .O(N__5175),
            .I(N__5160));
    LocalMux I__942 (
            .O(N__5172),
            .I(N__5157));
    InMux I__941 (
            .O(N__5171),
            .I(N__5154));
    LocalMux I__940 (
            .O(N__5168),
            .I(N__5149));
    LocalMux I__939 (
            .O(N__5165),
            .I(N__5149));
    Span4Mux_v I__938 (
            .O(N__5160),
            .I(N__5146));
    Span4Mux_h I__937 (
            .O(N__5157),
            .I(N__5143));
    LocalMux I__936 (
            .O(N__5154),
            .I(\uut.acc_out_1 ));
    Odrv12 I__935 (
            .O(N__5149),
            .I(\uut.acc_out_1 ));
    Odrv4 I__934 (
            .O(N__5146),
            .I(\uut.acc_out_1 ));
    Odrv4 I__933 (
            .O(N__5143),
            .I(\uut.acc_out_1 ));
    CascadeMux I__932 (
            .O(N__5134),
            .I(\uut.ALU_main.ALU_Out_0Z0Z_1_cascade_ ));
    InMux I__931 (
            .O(N__5131),
            .I(N__5128));
    LocalMux I__930 (
            .O(N__5128),
            .I(N__5125));
    Span4Mux_s2_h I__929 (
            .O(N__5125),
            .I(N__5121));
    InMux I__928 (
            .O(N__5124),
            .I(N__5118));
    Odrv4 I__927 (
            .O(N__5121),
            .I(\uut.un1_A_cry_0_c_RNI3CH45 ));
    LocalMux I__926 (
            .O(N__5118),
            .I(\uut.un1_A_cry_0_c_RNI3CH45 ));
    InMux I__925 (
            .O(N__5113),
            .I(N__5110));
    LocalMux I__924 (
            .O(N__5110),
            .I(N__5107));
    Span4Mux_v I__923 (
            .O(N__5107),
            .I(N__5104));
    Odrv4 I__922 (
            .O(N__5104),
            .I(\uut.seq.counter.un2_MAR_LD ));
    InMux I__921 (
            .O(N__5101),
            .I(N__5096));
    CascadeMux I__920 (
            .O(N__5100),
            .I(N__5093));
    InMux I__919 (
            .O(N__5099),
            .I(N__5089));
    LocalMux I__918 (
            .O(N__5096),
            .I(N__5086));
    InMux I__917 (
            .O(N__5093),
            .I(N__5083));
    CascadeMux I__916 (
            .O(N__5092),
            .I(N__5077));
    LocalMux I__915 (
            .O(N__5089),
            .I(N__5074));
    Span4Mux_v I__914 (
            .O(N__5086),
            .I(N__5069));
    LocalMux I__913 (
            .O(N__5083),
            .I(N__5069));
    InMux I__912 (
            .O(N__5082),
            .I(N__5064));
    InMux I__911 (
            .O(N__5081),
            .I(N__5064));
    InMux I__910 (
            .O(N__5080),
            .I(N__5061));
    InMux I__909 (
            .O(N__5077),
            .I(N__5058));
    Odrv12 I__908 (
            .O(N__5074),
            .I(\uut.T_2_rep1 ));
    Odrv4 I__907 (
            .O(N__5069),
            .I(\uut.T_2_rep1 ));
    LocalMux I__906 (
            .O(N__5064),
            .I(\uut.T_2_rep1 ));
    LocalMux I__905 (
            .O(N__5061),
            .I(\uut.T_2_rep1 ));
    LocalMux I__904 (
            .O(N__5058),
            .I(\uut.T_2_rep1 ));
    InMux I__903 (
            .O(N__5047),
            .I(N__5044));
    LocalMux I__902 (
            .O(N__5044),
            .I(\uut.seq.counter.T_2_rep1_RNIV9NUZ0 ));
    InMux I__901 (
            .O(N__5041),
            .I(N__5038));
    LocalMux I__900 (
            .O(N__5038),
            .I(N__5035));
    Span4Mux_h I__899 (
            .O(N__5035),
            .I(N__5032));
    Odrv4 I__898 (
            .O(N__5032),
            .I(\uut.bus_5 ));
    CascadeMux I__897 (
            .O(N__5029),
            .I(N__5025));
    CascadeMux I__896 (
            .O(N__5028),
            .I(N__5022));
    InMux I__895 (
            .O(N__5025),
            .I(N__5016));
    InMux I__894 (
            .O(N__5022),
            .I(N__5016));
    CascadeMux I__893 (
            .O(N__5021),
            .I(N__5013));
    LocalMux I__892 (
            .O(N__5016),
            .I(N__5009));
    InMux I__891 (
            .O(N__5013),
            .I(N__5006));
    InMux I__890 (
            .O(N__5012),
            .I(N__5003));
    Odrv4 I__889 (
            .O(N__5009),
            .I(\uut.q_0_fast_1 ));
    LocalMux I__888 (
            .O(N__5006),
            .I(\uut.q_0_fast_1 ));
    LocalMux I__887 (
            .O(N__5003),
            .I(\uut.q_0_fast_1 ));
    InMux I__886 (
            .O(N__4996),
            .I(N__4993));
    LocalMux I__885 (
            .O(N__4993),
            .I(\uut.seq.counter.T_1_fastZ0Z_0 ));
    InMux I__884 (
            .O(N__4990),
            .I(N__4983));
    InMux I__883 (
            .O(N__4989),
            .I(N__4983));
    CascadeMux I__882 (
            .O(N__4988),
            .I(N__4974));
    LocalMux I__881 (
            .O(N__4983),
            .I(N__4971));
    InMux I__880 (
            .O(N__4982),
            .I(N__4968));
    InMux I__879 (
            .O(N__4981),
            .I(N__4965));
    InMux I__878 (
            .O(N__4980),
            .I(N__4962));
    InMux I__877 (
            .O(N__4979),
            .I(N__4959));
    InMux I__876 (
            .O(N__4978),
            .I(N__4954));
    InMux I__875 (
            .O(N__4977),
            .I(N__4954));
    InMux I__874 (
            .O(N__4974),
            .I(N__4951));
    Odrv12 I__873 (
            .O(N__4971),
            .I(\uut.ir_out_fast_4 ));
    LocalMux I__872 (
            .O(N__4968),
            .I(\uut.ir_out_fast_4 ));
    LocalMux I__871 (
            .O(N__4965),
            .I(\uut.ir_out_fast_4 ));
    LocalMux I__870 (
            .O(N__4962),
            .I(\uut.ir_out_fast_4 ));
    LocalMux I__869 (
            .O(N__4959),
            .I(\uut.ir_out_fast_4 ));
    LocalMux I__868 (
            .O(N__4954),
            .I(\uut.ir_out_fast_4 ));
    LocalMux I__867 (
            .O(N__4951),
            .I(\uut.ir_out_fast_4 ));
    InMux I__866 (
            .O(N__4936),
            .I(N__4933));
    LocalMux I__865 (
            .O(N__4933),
            .I(N__4925));
    InMux I__864 (
            .O(N__4932),
            .I(N__4922));
    InMux I__863 (
            .O(N__4931),
            .I(N__4917));
    InMux I__862 (
            .O(N__4930),
            .I(N__4917));
    InMux I__861 (
            .O(N__4929),
            .I(N__4914));
    InMux I__860 (
            .O(N__4928),
            .I(N__4911));
    Span4Mux_h I__859 (
            .O(N__4925),
            .I(N__4901));
    LocalMux I__858 (
            .O(N__4922),
            .I(N__4901));
    LocalMux I__857 (
            .O(N__4917),
            .I(N__4898));
    LocalMux I__856 (
            .O(N__4914),
            .I(N__4893));
    LocalMux I__855 (
            .O(N__4911),
            .I(N__4893));
    InMux I__854 (
            .O(N__4910),
            .I(N__4888));
    InMux I__853 (
            .O(N__4909),
            .I(N__4888));
    InMux I__852 (
            .O(N__4908),
            .I(N__4881));
    InMux I__851 (
            .O(N__4907),
            .I(N__4881));
    InMux I__850 (
            .O(N__4906),
            .I(N__4881));
    Odrv4 I__849 (
            .O(N__4901),
            .I(\uut.ir_out_5 ));
    Odrv12 I__848 (
            .O(N__4898),
            .I(\uut.ir_out_5 ));
    Odrv4 I__847 (
            .O(N__4893),
            .I(\uut.ir_out_5 ));
    LocalMux I__846 (
            .O(N__4888),
            .I(\uut.ir_out_5 ));
    LocalMux I__845 (
            .O(N__4881),
            .I(\uut.ir_out_5 ));
    InMux I__844 (
            .O(N__4870),
            .I(N__4866));
    InMux I__843 (
            .O(N__4869),
            .I(N__4860));
    LocalMux I__842 (
            .O(N__4866),
            .I(N__4857));
    InMux I__841 (
            .O(N__4865),
            .I(N__4850));
    InMux I__840 (
            .O(N__4864),
            .I(N__4850));
    InMux I__839 (
            .O(N__4863),
            .I(N__4850));
    LocalMux I__838 (
            .O(N__4860),
            .I(\uut.q_ret_1_fast ));
    Odrv4 I__837 (
            .O(N__4857),
            .I(\uut.q_ret_1_fast ));
    LocalMux I__836 (
            .O(N__4850),
            .I(\uut.q_ret_1_fast ));
    InMux I__835 (
            .O(N__4843),
            .I(N__4836));
    InMux I__834 (
            .O(N__4842),
            .I(N__4833));
    InMux I__833 (
            .O(N__4841),
            .I(N__4830));
    InMux I__832 (
            .O(N__4840),
            .I(N__4827));
    InMux I__831 (
            .O(N__4839),
            .I(N__4824));
    LocalMux I__830 (
            .O(N__4836),
            .I(\uut.seq.counter.T_4 ));
    LocalMux I__829 (
            .O(N__4833),
            .I(\uut.seq.counter.T_4 ));
    LocalMux I__828 (
            .O(N__4830),
            .I(\uut.seq.counter.T_4 ));
    LocalMux I__827 (
            .O(N__4827),
            .I(\uut.seq.counter.T_4 ));
    LocalMux I__826 (
            .O(N__4824),
            .I(\uut.seq.counter.T_4 ));
    CascadeMux I__825 (
            .O(N__4813),
            .I(\uut.seq.un10_ACC_LD_xZ0Z1_cascade_ ));
    CascadeMux I__824 (
            .O(N__4810),
            .I(\uut.T_1_fast_RNI28LI1_0_cascade_ ));
    InMux I__823 (
            .O(N__4807),
            .I(N__4800));
    InMux I__822 (
            .O(N__4806),
            .I(N__4800));
    InMux I__821 (
            .O(N__4805),
            .I(N__4797));
    LocalMux I__820 (
            .O(N__4800),
            .I(N__4792));
    LocalMux I__819 (
            .O(N__4797),
            .I(N__4792));
    Span4Mux_v I__818 (
            .O(N__4792),
            .I(N__4789));
    Odrv4 I__817 (
            .O(N__4789),
            .I(\uut.N_41 ));
    CascadeMux I__816 (
            .O(N__4786),
            .I(\uut.seq.counter.T_2_rep1_RNIJDGJZ0_cascade_ ));
    InMux I__815 (
            .O(N__4783),
            .I(N__4779));
    InMux I__814 (
            .O(N__4782),
            .I(N__4776));
    LocalMux I__813 (
            .O(N__4779),
            .I(\uut.seq.D_4 ));
    LocalMux I__812 (
            .O(N__4776),
            .I(\uut.seq.D_4 ));
    CascadeMux I__811 (
            .O(N__4771),
            .I(\uut.D_1_3_cascade_ ));
    InMux I__810 (
            .O(N__4768),
            .I(N__4764));
    InMux I__809 (
            .O(N__4767),
            .I(N__4761));
    LocalMux I__808 (
            .O(N__4764),
            .I(N__4754));
    LocalMux I__807 (
            .O(N__4761),
            .I(N__4751));
    InMux I__806 (
            .O(N__4760),
            .I(N__4746));
    InMux I__805 (
            .O(N__4759),
            .I(N__4746));
    CascadeMux I__804 (
            .O(N__4758),
            .I(N__4743));
    CascadeMux I__803 (
            .O(N__4757),
            .I(N__4740));
    Span4Mux_h I__802 (
            .O(N__4754),
            .I(N__4733));
    Span4Mux_h I__801 (
            .O(N__4751),
            .I(N__4730));
    LocalMux I__800 (
            .O(N__4746),
            .I(N__4727));
    InMux I__799 (
            .O(N__4743),
            .I(N__4714));
    InMux I__798 (
            .O(N__4740),
            .I(N__4714));
    InMux I__797 (
            .O(N__4739),
            .I(N__4714));
    InMux I__796 (
            .O(N__4738),
            .I(N__4714));
    InMux I__795 (
            .O(N__4737),
            .I(N__4714));
    InMux I__794 (
            .O(N__4736),
            .I(N__4714));
    Odrv4 I__793 (
            .O(N__4733),
            .I(\uut.un7_ACC_LD ));
    Odrv4 I__792 (
            .O(N__4730),
            .I(\uut.un7_ACC_LD ));
    Odrv4 I__791 (
            .O(N__4727),
            .I(\uut.un7_ACC_LD ));
    LocalMux I__790 (
            .O(N__4714),
            .I(\uut.un7_ACC_LD ));
    InMux I__789 (
            .O(N__4705),
            .I(N__4697));
    InMux I__788 (
            .O(N__4704),
            .I(N__4692));
    InMux I__787 (
            .O(N__4703),
            .I(N__4692));
    InMux I__786 (
            .O(N__4702),
            .I(N__4689));
    InMux I__785 (
            .O(N__4701),
            .I(N__4686));
    InMux I__784 (
            .O(N__4700),
            .I(N__4681));
    LocalMux I__783 (
            .O(N__4697),
            .I(N__4678));
    LocalMux I__782 (
            .O(N__4692),
            .I(N__4674));
    LocalMux I__781 (
            .O(N__4689),
            .I(N__4671));
    LocalMux I__780 (
            .O(N__4686),
            .I(N__4668));
    InMux I__779 (
            .O(N__4685),
            .I(N__4663));
    InMux I__778 (
            .O(N__4684),
            .I(N__4663));
    LocalMux I__777 (
            .O(N__4681),
            .I(N__4658));
    Span4Mux_h I__776 (
            .O(N__4678),
            .I(N__4658));
    InMux I__775 (
            .O(N__4677),
            .I(N__4655));
    Odrv4 I__774 (
            .O(N__4674),
            .I(\uut.ir_out_4 ));
    Odrv4 I__773 (
            .O(N__4671),
            .I(\uut.ir_out_4 ));
    Odrv12 I__772 (
            .O(N__4668),
            .I(\uut.ir_out_4 ));
    LocalMux I__771 (
            .O(N__4663),
            .I(\uut.ir_out_4 ));
    Odrv4 I__770 (
            .O(N__4658),
            .I(\uut.ir_out_4 ));
    LocalMux I__769 (
            .O(N__4655),
            .I(\uut.ir_out_4 ));
    InMux I__768 (
            .O(N__4642),
            .I(N__4638));
    InMux I__767 (
            .O(N__4641),
            .I(N__4635));
    LocalMux I__766 (
            .O(N__4638),
            .I(\uut.seq.counter.T_1_fastZ0Z_3 ));
    LocalMux I__765 (
            .O(N__4635),
            .I(\uut.seq.counter.T_1_fastZ0Z_3 ));
    CascadeMux I__764 (
            .O(N__4630),
            .I(\uut.seq.counter.T_4_cascade_ ));
    InMux I__763 (
            .O(N__4627),
            .I(N__4624));
    LocalMux I__762 (
            .O(N__4624),
            .I(N__4621));
    Span4Mux_s3_h I__761 (
            .O(N__4621),
            .I(N__4618));
    Odrv4 I__760 (
            .O(N__4618),
            .I(\uut.seq.counter.T_1_fast_RNI4JTR1_0Z0Z_0 ));
    InMux I__759 (
            .O(N__4615),
            .I(N__4612));
    LocalMux I__758 (
            .O(N__4612),
            .I(N__4609));
    Span4Mux_h I__757 (
            .O(N__4609),
            .I(N__4606));
    Odrv4 I__756 (
            .O(N__4606),
            .I(\uut.ALU_main.un1_A_cry_5_c_RNINKZ0Z655 ));
    InMux I__755 (
            .O(N__4603),
            .I(\uut.ALU_main.un1_A_cry_5 ));
    InMux I__754 (
            .O(N__4600),
            .I(bfn_9_13_0_));
    InMux I__753 (
            .O(N__4597),
            .I(N__4594));
    LocalMux I__752 (
            .O(N__4594),
            .I(N__4591));
    Odrv12 I__751 (
            .O(N__4591),
            .I(\uut.ALU_main.un1_A_cry_6_c_RNINIMNZ0Z4 ));
    InMux I__750 (
            .O(N__4588),
            .I(N__4585));
    LocalMux I__749 (
            .O(N__4585),
            .I(\uut.ALU_main.un1_A_axb_1_l_ofxZ0 ));
    InMux I__748 (
            .O(N__4582),
            .I(N__4578));
    InMux I__747 (
            .O(N__4581),
            .I(N__4575));
    LocalMux I__746 (
            .O(N__4578),
            .I(N__4572));
    LocalMux I__745 (
            .O(N__4575),
            .I(N__4569));
    Odrv4 I__744 (
            .O(N__4572),
            .I(\uut.b_reg_out_6 ));
    Odrv12 I__743 (
            .O(N__4569),
            .I(\uut.b_reg_out_6 ));
    InMux I__742 (
            .O(N__4564),
            .I(N__4561));
    LocalMux I__741 (
            .O(N__4561),
            .I(\uut.ALU_main.un1_A_axb_6_l_ofxZ0 ));
    InMux I__740 (
            .O(N__4558),
            .I(N__4555));
    LocalMux I__739 (
            .O(N__4555),
            .I(N__4551));
    InMux I__738 (
            .O(N__4554),
            .I(N__4548));
    Span4Mux_h I__737 (
            .O(N__4551),
            .I(N__4545));
    LocalMux I__736 (
            .O(N__4548),
            .I(\uut.b_reg_out_5 ));
    Odrv4 I__735 (
            .O(N__4545),
            .I(\uut.b_reg_out_5 ));
    InMux I__734 (
            .O(N__4540),
            .I(N__4537));
    LocalMux I__733 (
            .O(N__4537),
            .I(\uut.ALU_main.un1_A_axb_5_l_ofxZ0 ));
    CascadeMux I__732 (
            .O(N__4534),
            .I(N__4531));
    InMux I__731 (
            .O(N__4531),
            .I(N__4528));
    LocalMux I__730 (
            .O(N__4528),
            .I(\uut.ALU_main.un1_A_axb_0_l_ofxZ0 ));
    InMux I__729 (
            .O(N__4525),
            .I(N__4521));
    InMux I__728 (
            .O(N__4524),
            .I(N__4518));
    LocalMux I__727 (
            .O(N__4521),
            .I(N__4515));
    LocalMux I__726 (
            .O(N__4518),
            .I(\uut.b_reg_out_7 ));
    Odrv12 I__725 (
            .O(N__4515),
            .I(\uut.b_reg_out_7 ));
    InMux I__724 (
            .O(N__4510),
            .I(N__4507));
    LocalMux I__723 (
            .O(N__4507),
            .I(\uut.ALU_main.un1_A_axbZ0Z_7 ));
    InMux I__722 (
            .O(N__4504),
            .I(N__4501));
    LocalMux I__721 (
            .O(N__4501),
            .I(N__4496));
    InMux I__720 (
            .O(N__4500),
            .I(N__4493));
    InMux I__719 (
            .O(N__4499),
            .I(N__4490));
    Span4Mux_h I__718 (
            .O(N__4496),
            .I(N__4487));
    LocalMux I__717 (
            .O(N__4493),
            .I(\uut.b_reg_out_2 ));
    LocalMux I__716 (
            .O(N__4490),
            .I(\uut.b_reg_out_2 ));
    Odrv4 I__715 (
            .O(N__4487),
            .I(\uut.b_reg_out_2 ));
    CascadeMux I__714 (
            .O(N__4480),
            .I(N__4475));
    CascadeMux I__713 (
            .O(N__4479),
            .I(N__4472));
    InMux I__712 (
            .O(N__4478),
            .I(N__4469));
    InMux I__711 (
            .O(N__4475),
            .I(N__4463));
    InMux I__710 (
            .O(N__4472),
            .I(N__4460));
    LocalMux I__709 (
            .O(N__4469),
            .I(N__4457));
    InMux I__708 (
            .O(N__4468),
            .I(N__4454));
    InMux I__707 (
            .O(N__4467),
            .I(N__4451));
    InMux I__706 (
            .O(N__4466),
            .I(N__4448));
    LocalMux I__705 (
            .O(N__4463),
            .I(N__4443));
    LocalMux I__704 (
            .O(N__4460),
            .I(N__4443));
    Span4Mux_v I__703 (
            .O(N__4457),
            .I(N__4438));
    LocalMux I__702 (
            .O(N__4454),
            .I(N__4438));
    LocalMux I__701 (
            .O(N__4451),
            .I(N__4435));
    LocalMux I__700 (
            .O(N__4448),
            .I(N__4430));
    Span4Mux_v I__699 (
            .O(N__4443),
            .I(N__4430));
    Odrv4 I__698 (
            .O(N__4438),
            .I(\uut.acc_out_2 ));
    Odrv4 I__697 (
            .O(N__4435),
            .I(\uut.acc_out_2 ));
    Odrv4 I__696 (
            .O(N__4430),
            .I(\uut.acc_out_2 ));
    InMux I__695 (
            .O(N__4423),
            .I(N__4420));
    LocalMux I__694 (
            .O(N__4420),
            .I(N__4412));
    InMux I__693 (
            .O(N__4419),
            .I(N__4409));
    InMux I__692 (
            .O(N__4418),
            .I(N__4406));
    InMux I__691 (
            .O(N__4417),
            .I(N__4401));
    InMux I__690 (
            .O(N__4416),
            .I(N__4401));
    CascadeMux I__689 (
            .O(N__4415),
            .I(N__4393));
    Span4Mux_v I__688 (
            .O(N__4412),
            .I(N__4390));
    LocalMux I__687 (
            .O(N__4409),
            .I(N__4385));
    LocalMux I__686 (
            .O(N__4406),
            .I(N__4385));
    LocalMux I__685 (
            .O(N__4401),
            .I(N__4382));
    InMux I__684 (
            .O(N__4400),
            .I(N__4371));
    InMux I__683 (
            .O(N__4399),
            .I(N__4371));
    InMux I__682 (
            .O(N__4398),
            .I(N__4371));
    InMux I__681 (
            .O(N__4397),
            .I(N__4371));
    InMux I__680 (
            .O(N__4396),
            .I(N__4371));
    InMux I__679 (
            .O(N__4393),
            .I(N__4368));
    Odrv4 I__678 (
            .O(N__4390),
            .I(\uut.un13_ACC_LD ));
    Odrv4 I__677 (
            .O(N__4385),
            .I(\uut.un13_ACC_LD ));
    Odrv4 I__676 (
            .O(N__4382),
            .I(\uut.un13_ACC_LD ));
    LocalMux I__675 (
            .O(N__4371),
            .I(\uut.un13_ACC_LD ));
    LocalMux I__674 (
            .O(N__4368),
            .I(\uut.un13_ACC_LD ));
    InMux I__673 (
            .O(N__4357),
            .I(N__4354));
    LocalMux I__672 (
            .O(N__4354),
            .I(\uut.ALU_main.un1_A_axb_2_l_ofxZ0 ));
    InMux I__671 (
            .O(N__4351),
            .I(N__4348));
    LocalMux I__670 (
            .O(N__4348),
            .I(\uut.pc.program_counter_0_1_1 ));
    CascadeMux I__669 (
            .O(N__4345),
            .I(N__4342));
    InMux I__668 (
            .O(N__4342),
            .I(N__4338));
    InMux I__667 (
            .O(N__4341),
            .I(N__4335));
    LocalMux I__666 (
            .O(N__4338),
            .I(N__4330));
    LocalMux I__665 (
            .O(N__4335),
            .I(N__4330));
    Odrv4 I__664 (
            .O(N__4330),
            .I(\uut.S0_0_i ));
    InMux I__663 (
            .O(N__4327),
            .I(N__4321));
    InMux I__662 (
            .O(N__4326),
            .I(N__4321));
    LocalMux I__661 (
            .O(N__4321),
            .I(N__4317));
    InMux I__660 (
            .O(N__4320),
            .I(N__4314));
    Odrv4 I__659 (
            .O(N__4317),
            .I(\uut.un1_A_cry_0_s ));
    LocalMux I__658 (
            .O(N__4314),
            .I(\uut.un1_A_cry_0_s ));
    InMux I__657 (
            .O(N__4309),
            .I(\uut.ALU_main.un1_A_cry_0_c_THRU_CO ));
    InMux I__656 (
            .O(N__4306),
            .I(\uut.ALU_main.un1_A_cry_0 ));
    InMux I__655 (
            .O(N__4303),
            .I(N__4300));
    LocalMux I__654 (
            .O(N__4300),
            .I(N__4297));
    Span4Mux_v I__653 (
            .O(N__4297),
            .I(N__4293));
    InMux I__652 (
            .O(N__4296),
            .I(N__4290));
    Odrv4 I__651 (
            .O(N__4293),
            .I(\uut.ALU_main.un1_A_cry_1_c_RNI7KLZ0Z45 ));
    LocalMux I__650 (
            .O(N__4290),
            .I(\uut.ALU_main.un1_A_cry_1_c_RNI7KLZ0Z45 ));
    InMux I__649 (
            .O(N__4285),
            .I(\uut.ALU_main.un1_A_cry_1 ));
    InMux I__648 (
            .O(N__4282),
            .I(N__4279));
    LocalMux I__647 (
            .O(N__4279),
            .I(\uut.ALU_main.un1_A_axb_3_l_ofxZ0 ));
    InMux I__646 (
            .O(N__4276),
            .I(\uut.ALU_main.un1_A_cry_2_cZ0 ));
    InMux I__645 (
            .O(N__4273),
            .I(N__4270));
    LocalMux I__644 (
            .O(N__4270),
            .I(N__4267));
    Odrv4 I__643 (
            .O(N__4267),
            .I(\uut.ALU_main.un1_A_axb_4_l_ofxZ0 ));
    InMux I__642 (
            .O(N__4264),
            .I(N__4261));
    LocalMux I__641 (
            .O(N__4261),
            .I(N__4258));
    Odrv4 I__640 (
            .O(N__4258),
            .I(\uut.ALU_main.un1_A_cry_3_c_RNIF4UZ0Z45 ));
    InMux I__639 (
            .O(N__4255),
            .I(\uut.ALU_main.un1_A_cry_3 ));
    InMux I__638 (
            .O(N__4252),
            .I(N__4249));
    LocalMux I__637 (
            .O(N__4249),
            .I(N__4246));
    Odrv4 I__636 (
            .O(N__4246),
            .I(\uut.ALU_main.un1_A_cry_4_c_RNIJCZ0Z255 ));
    InMux I__635 (
            .O(N__4243),
            .I(\uut.ALU_main.un1_A_cry_4 ));
    InMux I__634 (
            .O(N__4240),
            .I(N__4236));
    InMux I__633 (
            .O(N__4239),
            .I(N__4233));
    LocalMux I__632 (
            .O(N__4236),
            .I(N__4228));
    LocalMux I__631 (
            .O(N__4233),
            .I(N__4228));
    Odrv4 I__630 (
            .O(N__4228),
            .I(\uut.T_1_RNIVVKI3_3 ));
    InMux I__629 (
            .O(N__4225),
            .I(N__4220));
    InMux I__628 (
            .O(N__4224),
            .I(N__4215));
    InMux I__627 (
            .O(N__4223),
            .I(N__4215));
    LocalMux I__626 (
            .O(N__4220),
            .I(\uut.program_counter_m_0 ));
    LocalMux I__625 (
            .O(N__4215),
            .I(\uut.program_counter_m_0 ));
    CascadeMux I__624 (
            .O(N__4210),
            .I(\uut.pc.G_26_i_a4_5_sx_cascade_ ));
    InMux I__623 (
            .O(N__4207),
            .I(N__4204));
    LocalMux I__622 (
            .O(N__4204),
            .I(\uut.pc.G_26_i_a4_5 ));
    InMux I__621 (
            .O(N__4201),
            .I(N__4195));
    InMux I__620 (
            .O(N__4200),
            .I(N__4195));
    LocalMux I__619 (
            .O(N__4195),
            .I(N__4191));
    InMux I__618 (
            .O(N__4194),
            .I(N__4188));
    Odrv4 I__617 (
            .O(N__4191),
            .I(\uut.ir_out_m_c_c_0 ));
    LocalMux I__616 (
            .O(N__4188),
            .I(\uut.ir_out_m_c_c_0 ));
    InMux I__615 (
            .O(N__4183),
            .I(N__4180));
    LocalMux I__614 (
            .O(N__4180),
            .I(N__4177));
    Odrv4 I__613 (
            .O(N__4177),
            .I(\uut.alu_out_m_0_0 ));
    InMux I__612 (
            .O(N__4174),
            .I(N__4171));
    LocalMux I__611 (
            .O(N__4171),
            .I(N__4168));
    Span4Mux_h I__610 (
            .O(N__4168),
            .I(N__4165));
    Odrv4 I__609 (
            .O(N__4165),
            .I(\uut.alu_out_m_0 ));
    CascadeMux I__608 (
            .O(N__4162),
            .I(\uut.pc.program_counter_4_a1_0_0_1_cascade_ ));
    InMux I__607 (
            .O(N__4159),
            .I(N__4156));
    LocalMux I__606 (
            .O(N__4156),
            .I(\uut.pc.g2_0 ));
    InMux I__605 (
            .O(N__4153),
            .I(N__4150));
    LocalMux I__604 (
            .O(N__4150),
            .I(\uut.pc.N_77_0 ));
    CascadeMux I__603 (
            .O(N__4147),
            .I(\uut.pc.g1_0_cascade_ ));
    InMux I__602 (
            .O(N__4144),
            .I(N__4139));
    InMux I__601 (
            .O(N__4143),
            .I(N__4132));
    InMux I__600 (
            .O(N__4142),
            .I(N__4129));
    LocalMux I__599 (
            .O(N__4139),
            .I(N__4124));
    InMux I__598 (
            .O(N__4138),
            .I(N__4121));
    InMux I__597 (
            .O(N__4137),
            .I(N__4118));
    CascadeMux I__596 (
            .O(N__4136),
            .I(N__4113));
    InMux I__595 (
            .O(N__4135),
            .I(N__4110));
    LocalMux I__594 (
            .O(N__4132),
            .I(N__4107));
    LocalMux I__593 (
            .O(N__4129),
            .I(N__4104));
    CascadeMux I__592 (
            .O(N__4128),
            .I(N__4098));
    InMux I__591 (
            .O(N__4127),
            .I(N__4095));
    Span4Mux_h I__590 (
            .O(N__4124),
            .I(N__4092));
    LocalMux I__589 (
            .O(N__4121),
            .I(N__4087));
    LocalMux I__588 (
            .O(N__4118),
            .I(N__4087));
    InMux I__587 (
            .O(N__4117),
            .I(N__4080));
    InMux I__586 (
            .O(N__4116),
            .I(N__4080));
    InMux I__585 (
            .O(N__4113),
            .I(N__4080));
    LocalMux I__584 (
            .O(N__4110),
            .I(N__4073));
    Span4Mux_v I__583 (
            .O(N__4107),
            .I(N__4073));
    Span4Mux_v I__582 (
            .O(N__4104),
            .I(N__4073));
    InMux I__581 (
            .O(N__4103),
            .I(N__4070));
    InMux I__580 (
            .O(N__4102),
            .I(N__4067));
    InMux I__579 (
            .O(N__4101),
            .I(N__4062));
    InMux I__578 (
            .O(N__4098),
            .I(N__4062));
    LocalMux I__577 (
            .O(N__4095),
            .I(\uut.ir_out_7 ));
    Odrv4 I__576 (
            .O(N__4092),
            .I(\uut.ir_out_7 ));
    Odrv12 I__575 (
            .O(N__4087),
            .I(\uut.ir_out_7 ));
    LocalMux I__574 (
            .O(N__4080),
            .I(\uut.ir_out_7 ));
    Odrv4 I__573 (
            .O(N__4073),
            .I(\uut.ir_out_7 ));
    LocalMux I__572 (
            .O(N__4070),
            .I(\uut.ir_out_7 ));
    LocalMux I__571 (
            .O(N__4067),
            .I(\uut.ir_out_7 ));
    LocalMux I__570 (
            .O(N__4062),
            .I(\uut.ir_out_7 ));
    InMux I__569 (
            .O(N__4045),
            .I(N__4039));
    InMux I__568 (
            .O(N__4044),
            .I(N__4034));
    InMux I__567 (
            .O(N__4043),
            .I(N__4034));
    InMux I__566 (
            .O(N__4042),
            .I(N__4031));
    LocalMux I__565 (
            .O(N__4039),
            .I(N__4028));
    LocalMux I__564 (
            .O(N__4034),
            .I(N__4025));
    LocalMux I__563 (
            .O(N__4031),
            .I(N__4014));
    Span4Mux_h I__562 (
            .O(N__4028),
            .I(N__4014));
    Span4Mux_v I__561 (
            .O(N__4025),
            .I(N__4011));
    InMux I__560 (
            .O(N__4024),
            .I(N__4006));
    InMux I__559 (
            .O(N__4023),
            .I(N__4006));
    InMux I__558 (
            .O(N__4022),
            .I(N__4003));
    InMux I__557 (
            .O(N__4021),
            .I(N__3996));
    InMux I__556 (
            .O(N__4020),
            .I(N__3996));
    InMux I__555 (
            .O(N__4019),
            .I(N__3996));
    Odrv4 I__554 (
            .O(N__4014),
            .I(\uut.ir_out_6 ));
    Odrv4 I__553 (
            .O(N__4011),
            .I(\uut.ir_out_6 ));
    LocalMux I__552 (
            .O(N__4006),
            .I(\uut.ir_out_6 ));
    LocalMux I__551 (
            .O(N__4003),
            .I(\uut.ir_out_6 ));
    LocalMux I__550 (
            .O(N__3996),
            .I(\uut.ir_out_6 ));
    InMux I__549 (
            .O(N__3985),
            .I(N__3982));
    LocalMux I__548 (
            .O(N__3982),
            .I(\uut.AR_BUF.g0_3_a10_1Z0Z_1 ));
    InMux I__547 (
            .O(N__3979),
            .I(N__3975));
    InMux I__546 (
            .O(N__3978),
            .I(N__3972));
    LocalMux I__545 (
            .O(N__3975),
            .I(N__3969));
    LocalMux I__544 (
            .O(N__3972),
            .I(N__3966));
    Odrv12 I__543 (
            .O(N__3969),
            .I(\uut.D_1_0 ));
    Odrv4 I__542 (
            .O(N__3966),
            .I(\uut.D_1_0 ));
    CascadeMux I__541 (
            .O(N__3961),
            .I(\uut.AR_BUF.g0_3_a10_0Z0Z_2_cascade_ ));
    InMux I__540 (
            .O(N__3958),
            .I(N__3955));
    LocalMux I__539 (
            .O(N__3955),
            .I(\uut.AR_BUF.g0_3Z0Z_0 ));
    CascadeMux I__538 (
            .O(N__3952),
            .I(\uut.ir_out_m_c_d_0_cascade_ ));
    InMux I__537 (
            .O(N__3949),
            .I(N__3946));
    LocalMux I__536 (
            .O(N__3946),
            .I(\uut.AR_BUF.out_1_2_ivZ0Z_2 ));
    CascadeMux I__535 (
            .O(N__3943),
            .I(N__3940));
    InMux I__534 (
            .O(N__3940),
            .I(N__3937));
    LocalMux I__533 (
            .O(N__3937),
            .I(N__3934));
    Odrv4 I__532 (
            .O(N__3934),
            .I(\uut.AR_BUF.g0_1_a10_4Z0Z_1 ));
    CascadeMux I__531 (
            .O(N__3931),
            .I(\uut.AR_BUF.g0_3Z0Z_2_cascade_ ));
    CascadeMux I__530 (
            .O(N__3928),
            .I(\uut.AR_BUF.g0_3Z0Z_6_cascade_ ));
    InMux I__529 (
            .O(N__3925),
            .I(N__3920));
    InMux I__528 (
            .O(N__3924),
            .I(N__3915));
    InMux I__527 (
            .O(N__3923),
            .I(N__3915));
    LocalMux I__526 (
            .O(N__3920),
            .I(\uut.AR_out_0 ));
    LocalMux I__525 (
            .O(N__3915),
            .I(\uut.AR_out_0 ));
    CascadeMux I__524 (
            .O(N__3910),
            .I(\uut.seq.counter.un4_ACC_LD_cascade_ ));
    CascadeMux I__523 (
            .O(N__3907),
            .I(N__3904));
    InMux I__522 (
            .O(N__3904),
            .I(N__3901));
    LocalMux I__521 (
            .O(N__3901),
            .I(N__3898));
    Span4Mux_v I__520 (
            .O(N__3898),
            .I(N__3895));
    Odrv4 I__519 (
            .O(N__3895),
            .I(\uut.seq.counter.ACC_LD_0_0 ));
    InMux I__518 (
            .O(N__3892),
            .I(N__3888));
    InMux I__517 (
            .O(N__3891),
            .I(N__3885));
    LocalMux I__516 (
            .O(N__3888),
            .I(N__3880));
    LocalMux I__515 (
            .O(N__3885),
            .I(N__3877));
    InMux I__514 (
            .O(N__3884),
            .I(N__3874));
    InMux I__513 (
            .O(N__3883),
            .I(N__3871));
    Span4Mux_v I__512 (
            .O(N__3880),
            .I(N__3868));
    Span4Mux_h I__511 (
            .O(N__3877),
            .I(N__3863));
    LocalMux I__510 (
            .O(N__3874),
            .I(N__3863));
    LocalMux I__509 (
            .O(N__3871),
            .I(\uut.N_2_0 ));
    Odrv4 I__508 (
            .O(N__3868),
            .I(\uut.N_2_0 ));
    Odrv4 I__507 (
            .O(N__3863),
            .I(\uut.N_2_0 ));
    InMux I__506 (
            .O(N__3856),
            .I(N__3850));
    InMux I__505 (
            .O(N__3855),
            .I(N__3850));
    LocalMux I__504 (
            .O(N__3850),
            .I(N__3844));
    InMux I__503 (
            .O(N__3849),
            .I(N__3841));
    InMux I__502 (
            .O(N__3848),
            .I(N__3838));
    InMux I__501 (
            .O(N__3847),
            .I(N__3835));
    Odrv4 I__500 (
            .O(N__3844),
            .I(\uut.q_ret_1_fast_0 ));
    LocalMux I__499 (
            .O(N__3841),
            .I(\uut.q_ret_1_fast_0 ));
    LocalMux I__498 (
            .O(N__3838),
            .I(\uut.q_ret_1_fast_0 ));
    LocalMux I__497 (
            .O(N__3835),
            .I(\uut.q_ret_1_fast_0 ));
    CascadeMux I__496 (
            .O(N__3826),
            .I(\uut.AR_BUF.g0_3Z0Z_3_cascade_ ));
    InMux I__495 (
            .O(N__3823),
            .I(N__3820));
    LocalMux I__494 (
            .O(N__3820),
            .I(N__3817));
    Odrv4 I__493 (
            .O(N__3817),
            .I(\uut.AR_BUF.out_1_2_ivZ0Z_1 ));
    InMux I__492 (
            .O(N__3814),
            .I(N__3811));
    LocalMux I__491 (
            .O(N__3811),
            .I(N__3807));
    InMux I__490 (
            .O(N__3810),
            .I(N__3804));
    Span4Mux_v I__489 (
            .O(N__3807),
            .I(N__3798));
    LocalMux I__488 (
            .O(N__3804),
            .I(N__3798));
    CascadeMux I__487 (
            .O(N__3803),
            .I(N__3794));
    Span4Mux_v I__486 (
            .O(N__3798),
            .I(N__3791));
    InMux I__485 (
            .O(N__3797),
            .I(N__3788));
    InMux I__484 (
            .O(N__3794),
            .I(N__3785));
    Odrv4 I__483 (
            .O(N__3791),
            .I(\uut.un1_HLT_1 ));
    LocalMux I__482 (
            .O(N__3788),
            .I(\uut.un1_HLT_1 ));
    LocalMux I__481 (
            .O(N__3785),
            .I(\uut.un1_HLT_1 ));
    InMux I__480 (
            .O(N__3778),
            .I(N__3771));
    InMux I__479 (
            .O(N__3777),
            .I(N__3771));
    InMux I__478 (
            .O(N__3776),
            .I(N__3768));
    LocalMux I__477 (
            .O(N__3771),
            .I(N__3765));
    LocalMux I__476 (
            .O(N__3768),
            .I(\uut.N_5_0 ));
    Odrv4 I__475 (
            .O(N__3765),
            .I(\uut.N_5_0 ));
    InMux I__474 (
            .O(N__3760),
            .I(N__3757));
    LocalMux I__473 (
            .O(N__3757),
            .I(N__3754));
    Span4Mux_h I__472 (
            .O(N__3754),
            .I(N__3751));
    Odrv4 I__471 (
            .O(N__3751),
            .I(\uut.bus_6 ));
    InMux I__470 (
            .O(N__3748),
            .I(N__3745));
    LocalMux I__469 (
            .O(N__3745),
            .I(N__3742));
    Span4Mux_s2_v I__468 (
            .O(N__3742),
            .I(N__3739));
    Odrv4 I__467 (
            .O(N__3739),
            .I(\uut.bus_7 ));
    CascadeMux I__466 (
            .O(N__3736),
            .I(\uut.seq.D_2_0_x_cascade_ ));
    CascadeMux I__465 (
            .O(N__3733),
            .I(N__3728));
    CascadeMux I__464 (
            .O(N__3732),
            .I(N__3725));
    InMux I__463 (
            .O(N__3731),
            .I(N__3722));
    InMux I__462 (
            .O(N__3728),
            .I(N__3719));
    InMux I__461 (
            .O(N__3725),
            .I(N__3716));
    LocalMux I__460 (
            .O(N__3722),
            .I(\uut.q_0_fast ));
    LocalMux I__459 (
            .O(N__3719),
            .I(\uut.q_0_fast ));
    LocalMux I__458 (
            .O(N__3716),
            .I(\uut.q_0_fast ));
    InMux I__457 (
            .O(N__3709),
            .I(N__3703));
    InMux I__456 (
            .O(N__3708),
            .I(N__3703));
    LocalMux I__455 (
            .O(N__3703),
            .I(N__3700));
    Odrv4 I__454 (
            .O(N__3700),
            .I(\uut.data_1_2_ivdup ));
    CascadeMux I__453 (
            .O(N__3697),
            .I(\uut.IR.ir_out_m_c_d_1_3_cascade_ ));
    CascadeMux I__452 (
            .O(N__3694),
            .I(\uut.ir_out_m_c_d_3_cascade_ ));
    InMux I__451 (
            .O(N__3691),
            .I(N__3688));
    LocalMux I__450 (
            .O(N__3688),
            .I(\uut.seq.counter.T_2_rep1_RNIGC8CZ0Z1 ));
    CascadeMux I__449 (
            .O(N__3685),
            .I(\uut.seq.un13_ACC_LD_xZ0Z1_cascade_ ));
    CascadeMux I__448 (
            .O(N__3682),
            .I(\uut.seq.counter.T_2_rep1_RNI8TEZ0Z81_cascade_ ));
    CascadeMux I__447 (
            .O(N__3679),
            .I(\uut.seq.counter.un2_MAR_LD_cascade_ ));
    CascadeMux I__446 (
            .O(N__3676),
            .I(\uut.D_1_0_cascade_ ));
    InMux I__445 (
            .O(N__3673),
            .I(N__3670));
    LocalMux I__444 (
            .O(N__3670),
            .I(\uut.seq.q_ret_RNI52E81Z0Z_0 ));
    CascadeMux I__443 (
            .O(N__3667),
            .I(\uut.T_2_rep1_RNI6BLF1_cascade_ ));
    CascadeMux I__442 (
            .O(N__3664),
            .I(N__3661));
    InMux I__441 (
            .O(N__3661),
            .I(N__3658));
    LocalMux I__440 (
            .O(N__3658),
            .I(N__3655));
    Span4Mux_h I__439 (
            .O(N__3655),
            .I(N__3652));
    Odrv4 I__438 (
            .O(N__3652),
            .I(\uut.un17_IR_OE_0 ));
    InMux I__437 (
            .O(N__3649),
            .I(N__3645));
    CascadeMux I__436 (
            .O(N__3648),
            .I(N__3642));
    LocalMux I__435 (
            .O(N__3645),
            .I(N__3639));
    InMux I__434 (
            .O(N__3642),
            .I(N__3636));
    Odrv4 I__433 (
            .O(N__3639),
            .I(\uut.ir_out_m_d_0 ));
    LocalMux I__432 (
            .O(N__3636),
            .I(\uut.ir_out_m_d_0 ));
    CascadeMux I__431 (
            .O(N__3631),
            .I(\uut.pc.N_4_i_1_cascade_ ));
    InMux I__430 (
            .O(N__3628),
            .I(N__3624));
    InMux I__429 (
            .O(N__3627),
            .I(N__3621));
    LocalMux I__428 (
            .O(N__3624),
            .I(\uut.alu_out_m_2 ));
    LocalMux I__427 (
            .O(N__3621),
            .I(\uut.alu_out_m_2 ));
    CascadeMux I__426 (
            .O(N__3616),
            .I(\uut.ALU_main.N_43_0_cascade_ ));
    CascadeMux I__425 (
            .O(N__3613),
            .I(\uut.T_1_fast_RNIVM0N3_0_cascade_ ));
    InMux I__424 (
            .O(N__3610),
            .I(N__3607));
    LocalMux I__423 (
            .O(N__3607),
            .I(\uut.pc.N_11 ));
    CascadeMux I__422 (
            .O(N__3604),
            .I(\uut.AR_BUF.N_13_cascade_ ));
    CascadeMux I__421 (
            .O(N__3601),
            .I(\uut.AR_BUF.g0_1_0Z0Z_5_cascade_ ));
    InMux I__420 (
            .O(N__3598),
            .I(N__3595));
    LocalMux I__419 (
            .O(N__3595),
            .I(\uut.AR_BUF.g0_1_0Z0Z_1 ));
    CascadeMux I__418 (
            .O(N__3592),
            .I(N__3589));
    InMux I__417 (
            .O(N__3589),
            .I(N__3585));
    CascadeMux I__416 (
            .O(N__3588),
            .I(N__3581));
    LocalMux I__415 (
            .O(N__3585),
            .I(N__3578));
    InMux I__414 (
            .O(N__3584),
            .I(N__3573));
    InMux I__413 (
            .O(N__3581),
            .I(N__3573));
    Span4Mux_v I__412 (
            .O(N__3578),
            .I(N__3570));
    LocalMux I__411 (
            .O(N__3573),
            .I(\uut.AR_out_1 ));
    Odrv4 I__410 (
            .O(N__3570),
            .I(\uut.AR_out_1 ));
    InMux I__409 (
            .O(N__3565),
            .I(N__3562));
    LocalMux I__408 (
            .O(N__3562),
            .I(\uut.AR_BUF.g0_1_0_4_0 ));
    CascadeMux I__407 (
            .O(N__3559),
            .I(N__3554));
    CascadeMux I__406 (
            .O(N__3558),
            .I(N__3548));
    InMux I__405 (
            .O(N__3557),
            .I(N__3545));
    InMux I__404 (
            .O(N__3554),
            .I(N__3541));
    InMux I__403 (
            .O(N__3553),
            .I(N__3534));
    InMux I__402 (
            .O(N__3552),
            .I(N__3534));
    InMux I__401 (
            .O(N__3551),
            .I(N__3534));
    InMux I__400 (
            .O(N__3548),
            .I(N__3531));
    LocalMux I__399 (
            .O(N__3545),
            .I(N__3528));
    InMux I__398 (
            .O(N__3544),
            .I(N__3525));
    LocalMux I__397 (
            .O(N__3541),
            .I(N__3522));
    LocalMux I__396 (
            .O(N__3534),
            .I(N__3517));
    LocalMux I__395 (
            .O(N__3531),
            .I(N__3517));
    Sp12to4 I__394 (
            .O(N__3528),
            .I(N__3512));
    LocalMux I__393 (
            .O(N__3525),
            .I(N__3512));
    Span4Mux_v I__392 (
            .O(N__3522),
            .I(N__3507));
    Span4Mux_v I__391 (
            .O(N__3517),
            .I(N__3507));
    Odrv12 I__390 (
            .O(N__3512),
            .I(\uut.ir_out_1 ));
    Odrv4 I__389 (
            .O(N__3507),
            .I(\uut.ir_out_1 ));
    InMux I__388 (
            .O(N__3502),
            .I(N__3499));
    LocalMux I__387 (
            .O(N__3499),
            .I(\uut.AR_BUF.N_10 ));
    InMux I__386 (
            .O(N__3496),
            .I(N__3493));
    LocalMux I__385 (
            .O(N__3493),
            .I(\uut.AR_BUF.g0_1_0_0_0 ));
    InMux I__384 (
            .O(N__3490),
            .I(N__3487));
    LocalMux I__383 (
            .O(N__3487),
            .I(N__3484));
    Odrv4 I__382 (
            .O(N__3484),
            .I(\uut.AR_BUF.out_1_0_iv_2_1Z0Z_1 ));
    CascadeMux I__381 (
            .O(N__3481),
            .I(\uut.AR_BUF.g0_0_a5_0Z0Z_2_cascade_ ));
    InMux I__380 (
            .O(N__3478),
            .I(N__3475));
    LocalMux I__379 (
            .O(N__3475),
            .I(N__3472));
    Odrv12 I__378 (
            .O(N__3472),
            .I(\uut.AR_BUF.N_9 ));
    CascadeMux I__377 (
            .O(N__3469),
            .I(N__3466));
    InMux I__376 (
            .O(N__3466),
            .I(N__3463));
    LocalMux I__375 (
            .O(N__3463),
            .I(\uut.AR_BUF.g0_1_a10_3Z0Z_2 ));
    InMux I__374 (
            .O(N__3460),
            .I(N__3457));
    LocalMux I__373 (
            .O(N__3457),
            .I(\uut.AR_BUF.g0_0_o5_0Z0Z_0 ));
    CascadeMux I__372 (
            .O(N__3454),
            .I(\uut.AR_BUF.g0_1_a10_3_cascade_ ));
    InMux I__371 (
            .O(N__3451),
            .I(N__3448));
    LocalMux I__370 (
            .O(N__3448),
            .I(\uut.AR_BUF.N_7 ));
    InMux I__369 (
            .O(N__3445),
            .I(N__3439));
    InMux I__368 (
            .O(N__3444),
            .I(N__3439));
    LocalMux I__367 (
            .O(N__3439),
            .I(\uut.b_reg_out_4 ));
    InMux I__366 (
            .O(N__3436),
            .I(N__3433));
    LocalMux I__365 (
            .O(N__3433),
            .I(N__3430));
    Odrv12 I__364 (
            .O(N__3430),
            .I(\uut.AR_BUF.out_1_0_iv_2Z0Z_0 ));
    CascadeMux I__363 (
            .O(N__3427),
            .I(\uut.ir_out_m_d_2_cascade_ ));
    CascadeMux I__362 (
            .O(N__3424),
            .I(N__3421));
    InMux I__361 (
            .O(N__3421),
            .I(N__3418));
    LocalMux I__360 (
            .O(N__3418),
            .I(\uut.ALU_main.N_48 ));
    CascadeMux I__359 (
            .O(N__3415),
            .I(\uut.bus_6_cascade_ ));
    CascadeMux I__358 (
            .O(N__3412),
            .I(\uut.q_RNIDGA71_cascade_ ));
    CascadeMux I__357 (
            .O(N__3409),
            .I(\uut.ALU_main.N_45_cascade_ ));
    CascadeMux I__356 (
            .O(N__3406),
            .I(\uut.alu_out_m_4_cascade_ ));
    CascadeMux I__355 (
            .O(N__3403),
            .I(\uut.data_1_2_ivdup_cascade_ ));
    InMux I__354 (
            .O(N__3400),
            .I(N__3397));
    LocalMux I__353 (
            .O(N__3397),
            .I(\uut.N_4_0 ));
    InMux I__352 (
            .O(N__3394),
            .I(N__3391));
    LocalMux I__351 (
            .O(N__3391),
            .I(N__3388));
    Span4Mux_h I__350 (
            .O(N__3388),
            .I(N__3385));
    Odrv4 I__349 (
            .O(N__3385),
            .I(\uut.data_1_2_iv_0 ));
    CascadeMux I__348 (
            .O(N__3382),
            .I(\uut.program_counter_m_2_cascade_ ));
    InMux I__347 (
            .O(N__3379),
            .I(N__3376));
    LocalMux I__346 (
            .O(N__3376),
            .I(\uut.AR_BUF.N_8 ));
    CascadeMux I__345 (
            .O(N__3373),
            .I(N__3370));
    InMux I__344 (
            .O(N__3370),
            .I(N__3367));
    LocalMux I__343 (
            .O(N__3367),
            .I(\uut.program_counter_m_2 ));
    InMux I__342 (
            .O(N__3364),
            .I(N__3361));
    LocalMux I__341 (
            .O(N__3361),
            .I(\uut.AR_BUF.g0_0_0Z0Z_1 ));
    CascadeMux I__340 (
            .O(N__3358),
            .I(\uut.out_1_0_ivdup_2_cascade_ ));
    InMux I__339 (
            .O(N__3355),
            .I(N__3352));
    LocalMux I__338 (
            .O(N__3352),
            .I(\uut.ALU_main.N_43 ));
    InMux I__337 (
            .O(N__3349),
            .I(N__3346));
    LocalMux I__336 (
            .O(N__3346),
            .I(\uut.ir_out_m_d_1 ));
    CascadeMux I__335 (
            .O(N__3343),
            .I(\uut.acc_out_m_7_cascade_ ));
    CascadeMux I__334 (
            .O(N__3340),
            .I(\uut.bus_7_cascade_ ));
    InMux I__333 (
            .O(N__3337),
            .I(N__3334));
    LocalMux I__332 (
            .O(N__3334),
            .I(N__3331));
    Odrv4 I__331 (
            .O(N__3331),
            .I(\uut.N_1_0 ));
    IoInMux I__330 (
            .O(N__3328),
            .I(N__3325));
    LocalMux I__329 (
            .O(N__3325),
            .I(N__3322));
    Span4Mux_s2_h I__328 (
            .O(N__3322),
            .I(N__3319));
    Span4Mux_v I__327 (
            .O(N__3319),
            .I(N__3315));
    CascadeMux I__326 (
            .O(N__3318),
            .I(N__3312));
    Span4Mux_h I__325 (
            .O(N__3315),
            .I(N__3309));
    InMux I__324 (
            .O(N__3312),
            .I(N__3306));
    Odrv4 I__323 (
            .O(N__3309),
            .I(LED5_c));
    LocalMux I__322 (
            .O(N__3306),
            .I(LED5_c));
    CascadeMux I__321 (
            .O(N__3301),
            .I(\uut.out_1_2_iv_3_cascade_ ));
    IoInMux I__320 (
            .O(N__3298),
            .I(N__3295));
    LocalMux I__319 (
            .O(N__3295),
            .I(N__3292));
    Span4Mux_s2_h I__318 (
            .O(N__3292),
            .I(N__3289));
    Span4Mux_v I__317 (
            .O(N__3289),
            .I(N__3285));
    InMux I__316 (
            .O(N__3288),
            .I(N__3282));
    Odrv4 I__315 (
            .O(N__3285),
            .I(LED1_c));
    LocalMux I__314 (
            .O(N__3282),
            .I(LED1_c));
    CascadeMux I__313 (
            .O(N__3277),
            .I(\uut.ALU_main.N_47_cascade_ ));
    CascadeMux I__312 (
            .O(N__3274),
            .I(\uut.seq.un1_HLT_1_reti_cascade_ ));
    InMux I__311 (
            .O(N__3271),
            .I(N__3268));
    LocalMux I__310 (
            .O(N__3268),
            .I(N__3265));
    Odrv4 I__309 (
            .O(N__3265),
            .I(\uut.un1_HLT_0 ));
    CascadeMux I__308 (
            .O(N__3262),
            .I(\uut.ALU_main.N_46_cascade_ ));
    CascadeMux I__307 (
            .O(N__3259),
            .I(\uut.alu_out_m_5_cascade_ ));
    CascadeMux I__306 (
            .O(N__3256),
            .I(\uut.bus_5_cascade_ ));
    CascadeMux I__305 (
            .O(N__3253),
            .I(\uut.alu_out_m_7_cascade_ ));
    CascadeMux I__304 (
            .O(N__3250),
            .I(\uut.AR_BUF.out_1_1_iv_3_1Z0Z_0_cascade_ ));
    CascadeMux I__303 (
            .O(N__3247),
            .I(\uut.AR_BUF.out_1_1_ivZ0Z_0_cascade_ ));
    CascadeMux I__302 (
            .O(N__3244),
            .I(\uut.out_1_1_iv_2_cascade_ ));
    InMux I__301 (
            .O(N__3241),
            .I(N__3238));
    LocalMux I__300 (
            .O(N__3238),
            .I(G_138));
    CascadeMux I__299 (
            .O(N__3235),
            .I(G_138_cascade_));
    IoInMux I__298 (
            .O(N__3232),
            .I(N__3229));
    LocalMux I__297 (
            .O(N__3229),
            .I(N__3226));
    Odrv12 I__296 (
            .O(N__3226),
            .I(\uut.buf_clk_1 ));
    INV \INVuut.mar.ff4.q_neC  (
            .O(\INVuut.mar.ff4.q_neC_net ),
            .I(N__5658));
    INV \INVuut.out_reg.ff4.qC  (
            .O(\INVuut.out_reg.ff4.qC_net ),
            .I(N__5656));
    INV \INVuut.seq.counter.T_1_0C  (
            .O(\INVuut.seq.counter.T_1_0C_net ),
            .I(N__5652));
    INV \INVuut.AR.ff4.q_neC  (
            .O(\INVuut.AR.ff4.q_neC_net ),
            .I(N__5649));
    INV \INVuut.AR.ff3.qC  (
            .O(\INVuut.AR.ff3.qC_net ),
            .I(N__5645));
    INV \INVuut.IR.ff3.qC  (
            .O(\INVuut.IR.ff3.qC_net ),
            .I(N__5659));
    INV \INVuut.b_reg.ff1.qC  (
            .O(\INVuut.b_reg.ff1.qC_net ),
            .I(N__5657));
    INV \INVuut.out_reg.ff3.qC  (
            .O(\INVuut.out_reg.ff3.qC_net ),
            .I(N__5655));
    INV \INVuut.acc.ff4.qC  (
            .O(\INVuut.acc.ff4.qC_net ),
            .I(N__5651));
    INV \INVuut.mar.ff2.q_neC  (
            .O(\INVuut.mar.ff2.q_neC_net ),
            .I(N__5644));
    INV \INVuut.seq.counter.T_1_1C  (
            .O(\INVuut.seq.counter.T_1_1C_net ),
            .I(N__5641));
    INV \INVuut.seq.counter.T_1_4C  (
            .O(\INVuut.seq.counter.T_1_4C_net ),
            .I(N__5637));
    INV \INVuut.IR.ff6.q_0_fastC  (
            .O(\INVuut.IR.ff6.q_0_fastC_net ),
            .I(N__5654));
    INV \INVuut.b_reg.ff4.qC  (
            .O(\INVuut.b_reg.ff4.qC_net ),
            .I(N__5640));
    INV \INVuut.AR.ff1.q_neC  (
            .O(\INVuut.AR.ff1.q_neC_net ),
            .I(N__5635));
    INV \INVuut.acc.ff1.qC  (
            .O(\INVuut.acc.ff1.qC_net ),
            .I(N__5636));
    INV \INVuut.seq.counter.T_1_fast_3C  (
            .O(\INVuut.seq.counter.T_1_fast_3C_net ),
            .I(N__5653));
    INV \INVuut.IR.ff5.q_0_rep1C  (
            .O(\INVuut.IR.ff5.q_0_rep1C_net ),
            .I(N__5650));
    INV \INVuut.IR.ff7.q_ret_1_fastC  (
            .O(\INVuut.IR.ff7.q_ret_1_fastC_net ),
            .I(N__5647));
    INV \INVuut.IR.ff4.q_neC  (
            .O(\INVuut.IR.ff4.q_neC_net ),
            .I(N__5643));
    INV \INVuut.b_reg.ff3.qC  (
            .O(\INVuut.b_reg.ff3.qC_net ),
            .I(N__5634));
    INV \INVuut.IR.ff1.q_neC  (
            .O(\INVuut.IR.ff1.q_neC_net ),
            .I(N__5646));
    INV \INVuut.seq.q_retC  (
            .O(\INVuut.seq.q_retC_net ),
            .I(N__5642));
    INV \INVuut.IR.ff5.q_0_neC  (
            .O(\INVuut.IR.ff5.q_0_neC_net ),
            .I(N__5639));
    INV \INVuut.b_reg.ff5.qC  (
            .O(\INVuut.b_reg.ff5.qC_net ),
            .I(N__5633));
    INV \INVuut.acc.ff3.qC  (
            .O(\INVuut.acc.ff3.qC_net ),
            .I(N__5624));
    INV \INVuut.out_reg.ff1.qC  (
            .O(\INVuut.out_reg.ff1.qC_net ),
            .I(N__5628));
    INV \INVuut.out_reg.ff5.qC  (
            .O(\INVuut.out_reg.ff5.qC_net ),
            .I(N__5638));
    INV \INVuut.b_reg.ff8.qC  (
            .O(\INVuut.b_reg.ff8.qC_net ),
            .I(N__5632));
    INV \INVuut.seq.q_ret_1C  (
            .O(\INVuut.seq.q_ret_1C_net ),
            .I(N__5630));
    INV \INVuut.AR.ff2.qC  (
            .O(\INVuut.AR.ff2.qC_net ),
            .I(N__5625));
    INV \INVuut.acc.ff2.qC  (
            .O(\INVuut.acc.ff2.qC_net ),
            .I(N__5623));
    INV \INVuut.b_reg.ff7.qC  (
            .O(\INVuut.b_reg.ff7.qC_net ),
            .I(N__5629));
    INV \INVuut.b_reg.ff6.qC  (
            .O(\INVuut.b_reg.ff6.qC_net ),
            .I(N__5626));
    defparam IN_MUX_bfv_9_12_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_12_0_ (
            .carryinitin(),
            .carryinitout(bfn_9_12_0_));
    defparam IN_MUX_bfv_9_13_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_9_13_0_ (
            .carryinitin(\uut.ALU_main.un1_A_cry_6 ),
            .carryinitout(bfn_9_13_0_));
    ICE_GB \uut.buf_clk_1_inferred_clock_0_RNIQBSF  (
            .USERSIGNALTOGLOBALBUFFER(N__3232),
            .GLOBALBUFFEROUTPUT(\uut.buf_clk_1_g ));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam N_62_i_LC_5_9_1.C_ON=1'b0;
    defparam N_62_i_LC_5_9_1.SEQ_MODE=4'b0000;
    defparam N_62_i_LC_5_9_1.LUT_INIT=16'b0101010101010101;
    LogicCell40 N_62_i_LC_5_9_1 (
            .in0(N__3241),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(G_138),
            .ltout(G_138_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.buf_clk_1_inferred_clock_0_RNO_LC_5_9_2 .C_ON=1'b0;
    defparam \uut.buf_clk_1_inferred_clock_0_RNO_LC_5_9_2 .SEQ_MODE=4'b0000;
    defparam \uut.buf_clk_1_inferred_clock_0_RNO_LC_5_9_2 .LUT_INIT=16'b0101000001010000;
    LogicCell40 \uut.buf_clk_1_inferred_clock_0_RNO_LC_5_9_2  (
            .in0(N__3271),
            .in1(_gnd_net_),
            .in2(N__3235),
            .in3(_gnd_net_),
            .lcout(\uut.buf_clk_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.b_reg.ff6.q_LC_5_12_1 .C_ON=1'b0;
    defparam \uut.b_reg.ff6.q_LC_5_12_1 .SEQ_MODE=4'b1000;
    defparam \uut.b_reg.ff6.q_LC_5_12_1 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \uut.b_reg.ff6.q_LC_5_12_1  (
            .in0(N__6101),
            .in1(N__6128),
            .in2(N__6079),
            .in3(N__9044),
            .lcout(\uut.b_reg_out_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.b_reg.ff6.qC_net ),
            .ce(N__7515),
            .sr(_gnd_net_));
    defparam \uut.b_reg.ff7.q_LC_5_13_1 .C_ON=1'b0;
    defparam \uut.b_reg.ff7.q_LC_5_13_1 .SEQ_MODE=4'b1000;
    defparam \uut.b_reg.ff7.q_LC_5_13_1 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \uut.b_reg.ff7.q_LC_5_13_1  (
            .in0(N__6363),
            .in1(N__6402),
            .in2(N__6331),
            .in3(N__9045),
            .lcout(\uut.b_reg_out_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.b_reg.ff7.qC_net ),
            .ce(N__7514),
            .sr(_gnd_net_));
    defparam \uut.acc.ff2.q_LC_6_9_0 .C_ON=1'b0;
    defparam \uut.acc.ff2.q_LC_6_9_0 .SEQ_MODE=4'b1000;
    defparam \uut.acc.ff2.q_LC_6_9_0 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \uut.acc.ff2.q_LC_6_9_0  (
            .in0(N__7684),
            .in1(N__7644),
            .in2(_gnd_net_),
            .in3(N__7579),
            .lcout(\uut.acc_out_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.acc.ff2.qC_net ),
            .ce(N__5833),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.out_1_1_iv_3_1_0_LC_6_10_2 .C_ON=1'b0;
    defparam \uut.AR_BUF.out_1_1_iv_3_1_0_LC_6_10_2 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.out_1_1_iv_3_1_0_LC_6_10_2 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \uut.AR_BUF.out_1_1_iv_3_1_0_LC_6_10_2  (
            .in0(N__5171),
            .in1(N__8282),
            .in2(N__3588),
            .in3(N__7783),
            .lcout(),
            .ltout(\uut.AR_BUF.out_1_1_iv_3_1Z0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.out_1_1_iv_0_LC_6_10_3 .C_ON=1'b0;
    defparam \uut.AR_BUF.out_1_1_iv_0_LC_6_10_3 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.out_1_1_iv_0_LC_6_10_3 .LUT_INIT=16'b1111101111111010;
    LogicCell40 \uut.AR_BUF.out_1_1_iv_0_LC_6_10_3  (
            .in0(N__5750),
            .in1(N__7102),
            .in2(N__3250),
            .in3(N__3557),
            .lcout(),
            .ltout(\uut.AR_BUF.out_1_1_ivZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.out_1_1_iv_2_LC_6_10_4 .C_ON=1'b0;
    defparam \uut.AR_BUF.out_1_1_iv_2_LC_6_10_4 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.out_1_1_iv_2_LC_6_10_4 .LUT_INIT=16'b1111111111110001;
    LogicCell40 \uut.AR_BUF.out_1_1_iv_2_LC_6_10_4  (
            .in0(N__9072),
            .in1(N__6817),
            .in2(N__3247),
            .in3(N__3349),
            .lcout(),
            .ltout(\uut.out_1_1_iv_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR.ff2.q_LC_6_10_5 .C_ON=1'b0;
    defparam \uut.AR.ff2.q_LC_6_10_5 .SEQ_MODE=4'b1000;
    defparam \uut.AR.ff2.q_LC_6_10_5 .LUT_INIT=16'b1111101111001000;
    LogicCell40 \uut.AR.ff2.q_LC_6_10_5  (
            .in0(N__7692),
            .in1(N__8032),
            .in2(N__3244),
            .in3(N__3584),
            .lcout(\uut.AR_out_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.AR.ff2.qC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.acc.ff6.q_RNIEIB71_LC_6_11_2 .C_ON=1'b0;
    defparam \uut.acc.ff6.q_RNIEIB71_LC_6_11_2 .SEQ_MODE=4'b0000;
    defparam \uut.acc.ff6.q_RNIEIB71_LC_6_11_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uut.acc.ff6.q_RNIEIB71_LC_6_11_2  (
            .in0(N__6030),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8281),
            .lcout(\uut.acc_out_m_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.ALU_Out_0_6_LC_6_11_3 .C_ON=1'b0;
    defparam \uut.ALU_main.ALU_Out_0_6_LC_6_11_3 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.ALU_Out_0_6_LC_6_11_3 .LUT_INIT=16'b1000100001100110;
    LogicCell40 \uut.ALU_main.ALU_Out_0_6_LC_6_11_3  (
            .in0(N__6272),
            .in1(N__4582),
            .in2(_gnd_net_),
            .in3(N__6774),
            .lcout(),
            .ltout(\uut.ALU_main.N_47_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_cry_5_c_RNISM3EE_LC_6_11_4 .C_ON=1'b0;
    defparam \uut.ALU_main.un1_A_cry_5_c_RNISM3EE_LC_6_11_4 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_cry_5_c_RNISM3EE_LC_6_11_4 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \uut.ALU_main.un1_A_cry_5_c_RNISM3EE_LC_6_11_4  (
            .in0(N__4615),
            .in1(N__6616),
            .in2(N__3277),
            .in3(N__6492),
            .lcout(\uut.alu_out_m_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_RNIT9ANK_1_LC_6_12_1 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_RNIT9ANK_1_LC_6_12_1 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_RNIT9ANK_1_LC_6_12_1 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \uut.seq.counter.T_1_RNIT9ANK_1_LC_6_12_1  (
            .in0(_gnd_net_),
            .in1(N__7414),
            .in2(_gnd_net_),
            .in3(N__3883),
            .lcout(),
            .ltout(\uut.seq.un1_HLT_1_reti_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.q_ret_1_LC_6_12_2 .C_ON=1'b0;
    defparam \uut.seq.q_ret_1_LC_6_12_2 .SEQ_MODE=4'b1000;
    defparam \uut.seq.q_ret_1_LC_6_12_2 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uut.seq.q_ret_1_LC_6_12_2  (
            .in0(N__3776),
            .in1(N__3400),
            .in2(N__3274),
            .in3(N__3337),
            .lcout(\uut.un1_HLT_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.seq.q_ret_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.ALU_Out_0_5_LC_6_12_4 .C_ON=1'b0;
    defparam \uut.ALU_main.ALU_Out_0_5_LC_6_12_4 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.ALU_Out_0_5_LC_6_12_4 .LUT_INIT=16'b1000100001100110;
    LogicCell40 \uut.ALU_main.ALU_Out_0_5_LC_6_12_4  (
            .in0(N__4554),
            .in1(N__6029),
            .in2(_gnd_net_),
            .in3(N__6766),
            .lcout(),
            .ltout(\uut.ALU_main.N_46_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_cry_4_c_RNIMATDE_LC_6_12_5 .C_ON=1'b0;
    defparam \uut.ALU_main.un1_A_cry_4_c_RNIMATDE_LC_6_12_5 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_cry_4_c_RNIMATDE_LC_6_12_5 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \uut.ALU_main.un1_A_cry_4_c_RNIMATDE_LC_6_12_5  (
            .in0(N__4252),
            .in1(N__6620),
            .in2(N__3262),
            .in3(N__6502),
            .lcout(\uut.alu_out_m_5 ),
            .ltout(\uut.alu_out_m_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mem.data_1_1_iv_LC_6_12_6 .C_ON=1'b0;
    defparam \uut.mem.data_1_1_iv_LC_6_12_6 .SEQ_MODE=4'b0000;
    defparam \uut.mem.data_1_1_iv_LC_6_12_6 .LUT_INIT=16'b1111110011111101;
    LogicCell40 \uut.mem.data_1_1_iv_LC_6_12_6  (
            .in0(N__6074),
            .in1(N__6100),
            .in2(N__3259),
            .in3(N__9038),
            .lcout(\uut.bus_5 ),
            .ltout(\uut.bus_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff6.q_0_ne_RNIV8OLK_LC_6_12_7 .C_ON=1'b0;
    defparam \uut.IR.ff6.q_0_ne_RNIV8OLK_LC_6_12_7 .SEQ_MODE=4'b0000;
    defparam \uut.IR.ff6.q_0_ne_RNIV8OLK_LC_6_12_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \uut.IR.ff6.q_0_ne_RNIV8OLK_LC_6_12_7  (
            .in0(_gnd_net_),
            .in1(N__7413),
            .in2(N__3256),
            .in3(N__4936),
            .lcout(\uut.N_2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_cry_6_c_RNIUOL0E_LC_6_13_0 .C_ON=1'b0;
    defparam \uut.ALU_main.un1_A_cry_6_c_RNIUOL0E_LC_6_13_0 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_cry_6_c_RNIUOL0E_LC_6_13_0 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \uut.ALU_main.un1_A_cry_6_c_RNIUOL0E_LC_6_13_0  (
            .in0(N__4597),
            .in1(N__6619),
            .in2(N__3424),
            .in3(N__6501),
            .lcout(\uut.alu_out_m_7 ),
            .ltout(\uut.alu_out_m_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.b_reg.ff8.q_LC_6_13_1 .C_ON=1'b0;
    defparam \uut.b_reg.ff8.q_LC_6_13_1 .SEQ_MODE=4'b1000;
    defparam \uut.b_reg.ff8.q_LC_6_13_1 .LUT_INIT=16'b1111101011111011;
    LogicCell40 \uut.b_reg.ff8.q_LC_6_13_1  (
            .in0(N__6215),
            .in1(N__6889),
            .in2(N__3253),
            .in3(N__9074),
            .lcout(\uut.b_reg_out_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.b_reg.ff8.qC_net ),
            .ce(N__7503),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_RNI5ENL7_3_LC_6_13_7 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_RNI5ENL7_3_LC_6_13_7 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_RNI5ENL7_3_LC_6_13_7 .LUT_INIT=16'b1111111111101111;
    LogicCell40 \uut.seq.counter.T_1_RNI5ENL7_3_LC_6_13_7  (
            .in0(N__6760),
            .in1(N__4768),
            .in2(N__3907),
            .in3(N__4423),
            .lcout(\uut.ACC_LD_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.acc.ff8.q_RNIGMD71_LC_6_14_2 .C_ON=1'b0;
    defparam \uut.acc.ff8.q_RNIGMD71_LC_6_14_2 .SEQ_MODE=4'b0000;
    defparam \uut.acc.ff8.q_RNIGMD71_LC_6_14_2 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uut.acc.ff8.q_RNIGMD71_LC_6_14_2  (
            .in0(N__6178),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8273),
            .lcout(\uut.acc_out_m_7 ),
            .ltout(\uut.acc_out_m_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mem.data_1_iv_LC_6_14_3 .C_ON=1'b0;
    defparam \uut.mem.data_1_iv_LC_6_14_3 .SEQ_MODE=4'b0000;
    defparam \uut.mem.data_1_iv_LC_6_14_3 .LUT_INIT=16'b1111110011111101;
    LogicCell40 \uut.mem.data_1_iv_LC_6_14_3  (
            .in0(N__9005),
            .in1(N__6194),
            .in2(N__3343),
            .in3(N__6874),
            .lcout(\uut.bus_7 ),
            .ltout(\uut.bus_7_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff8.q_0_ne_RNIB9TFK_LC_6_14_4 .C_ON=1'b0;
    defparam \uut.IR.ff8.q_0_ne_RNIB9TFK_LC_6_14_4 .SEQ_MODE=4'b0000;
    defparam \uut.IR.ff8.q_0_ne_RNIB9TFK_LC_6_14_4 .LUT_INIT=16'b1111000011001100;
    LogicCell40 \uut.IR.ff8.q_0_ne_RNIB9TFK_LC_6_14_4  (
            .in0(_gnd_net_),
            .in1(N__4127),
            .in2(N__3340),
            .in3(N__7415),
            .lcout(\uut.N_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.out_reg.ff5.q_LC_6_14_7 .C_ON=1'b0;
    defparam \uut.out_reg.ff5.q_LC_6_14_7 .SEQ_MODE=4'b1000;
    defparam \uut.out_reg.ff5.q_LC_6_14_7 .LUT_INIT=16'b1111101011011000;
    LogicCell40 \uut.out_reg.ff5.q_LC_6_14_7  (
            .in0(N__8274),
            .in1(N__3394),
            .in2(N__3318),
            .in3(N__5913),
            .lcout(LED5_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.out_reg.ff5.qC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_1_a10_3_2_LC_7_8_2 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_1_a10_3_2_LC_7_8_2 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_1_a10_3_2_LC_7_8_2 .LUT_INIT=16'b0000000010001000;
    LogicCell40 \uut.AR_BUF.g0_1_a10_3_2_LC_7_8_2  (
            .in0(N__4701),
            .in1(N__3544),
            .in2(_gnd_net_),
            .in3(N__4137),
            .lcout(\uut.AR_BUF.g0_1_a10_3Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.out_1_2_iv_3_LC_7_8_6 .C_ON=1'b0;
    defparam \uut.AR_BUF.out_1_2_iv_3_LC_7_8_6 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.out_1_2_iv_3_LC_7_8_6 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \uut.AR_BUF.out_1_2_iv_3_LC_7_8_6  (
            .in0(N__4174),
            .in1(N__3823),
            .in2(_gnd_net_),
            .in3(N__3649),
            .lcout(),
            .ltout(\uut.out_1_2_iv_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.out_reg.ff1.q_LC_7_8_7 .C_ON=1'b0;
    defparam \uut.out_reg.ff1.q_LC_7_8_7 .SEQ_MODE=4'b1000;
    defparam \uut.out_reg.ff1.q_LC_7_8_7 .LUT_INIT=16'b1110111011100010;
    LogicCell40 \uut.out_reg.ff1.q_LC_7_8_7  (
            .in0(N__3288),
            .in1(N__8287),
            .in2(N__3301),
            .in3(N__9262),
            .lcout(LED1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.out_reg.ff1.qC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.acc.ff3.q_LC_7_9_1 .C_ON=1'b0;
    defparam \uut.acc.ff3.q_LC_7_9_1 .SEQ_MODE=4'b1000;
    defparam \uut.acc.ff3.q_LC_7_9_1 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \uut.acc.ff3.q_LC_7_9_1  (
            .in0(N__8098),
            .in1(N__3627),
            .in2(N__5452),
            .in3(N__9073),
            .lcout(\uut.acc_out_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.acc.ff3.qC_net ),
            .ce(N__5845),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_0_0_1_LC_7_9_2 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_0_0_1_LC_7_9_2 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_0_0_1_LC_7_9_2 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \uut.AR_BUF.g0_0_0_1_LC_7_9_2  (
            .in0(N__7762),
            .in1(N__4466),
            .in2(N__7171),
            .in3(N__8260),
            .lcout(\uut.AR_BUF.g0_0_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_0_a5_LC_7_9_4 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_0_a5_LC_7_9_4 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_0_a5_LC_7_9_4 .LUT_INIT=16'b1111000011100000;
    LogicCell40 \uut.AR_BUF.g0_0_a5_LC_7_9_4  (
            .in0(N__7974),
            .in1(N__3460),
            .in2(N__7258),
            .in3(N__8385),
            .lcout(\uut.AR_BUF.N_8 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_RNIEETC1_0_LC_7_10_0 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_RNIEETC1_0_LC_7_10_0 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_RNIEETC1_0_LC_7_10_0 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \uut.seq.counter.T_1_RNIEETC1_0_LC_7_10_0  (
            .in0(N__8756),
            .in1(N__8659),
            .in2(N__5792),
            .in3(N__8579),
            .lcout(\uut.program_counter_m_2 ),
            .ltout(\uut.program_counter_m_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.out_1_0_iv_2_0_LC_7_10_1 .C_ON=1'b0;
    defparam \uut.AR_BUF.out_1_0_iv_2_0_LC_7_10_1 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.out_1_0_iv_2_0_LC_7_10_1 .LUT_INIT=16'b1111110011110000;
    LogicCell40 \uut.AR_BUF.out_1_0_iv_2_0_LC_7_10_1  (
            .in0(_gnd_net_),
            .in1(N__7167),
            .in2(N__3382),
            .in3(N__7764),
            .lcout(\uut.AR_BUF.out_1_0_iv_2Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_cry_1_c_RNI46ADE_0_LC_7_10_2 .C_ON=1'b0;
    defparam \uut.ALU_main.un1_A_cry_1_c_RNI46ADE_0_LC_7_10_2 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_cry_1_c_RNI46ADE_0_LC_7_10_2 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \uut.ALU_main.un1_A_cry_1_c_RNI46ADE_0_LC_7_10_2  (
            .in0(N__6618),
            .in1(N__3355),
            .in2(N__6496),
            .in3(N__4303),
            .lcout(\uut.alu_out_m_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_0_0_LC_7_10_6 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_0_0_LC_7_10_6 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_0_0_LC_7_10_6 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uut.AR_BUF.g0_0_0_LC_7_10_6  (
            .in0(N__3379),
            .in1(N__3478),
            .in2(N__3373),
            .in3(N__3364),
            .lcout(\uut.out_1_0_ivdup_2 ),
            .ltout(\uut.out_1_0_ivdup_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.pc.program_counter_2_LC_7_10_7 .C_ON=1'b0;
    defparam \uut.pc.program_counter_2_LC_7_10_7 .SEQ_MODE=4'b1000;
    defparam \uut.pc.program_counter_2_LC_7_10_7 .LUT_INIT=16'b1011101110111001;
    LogicCell40 \uut.pc.program_counter_2_LC_7_10_7  (
            .in0(N__5485),
            .in1(N__5461),
            .in2(N__3358),
            .in3(N__7185),
            .lcout(\uut.program_counter_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5627),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.ALU_Out_0_2_LC_7_11_0 .C_ON=1'b0;
    defparam \uut.ALU_main.ALU_Out_0_2_LC_7_11_0 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.ALU_Out_0_2_LC_7_11_0 .LUT_INIT=16'b1000100001100110;
    LogicCell40 \uut.ALU_main.ALU_Out_0_2_LC_7_11_0  (
            .in0(N__4468),
            .in1(N__4500),
            .in2(_gnd_net_),
            .in3(N__6775),
            .lcout(\uut.ALU_main.N_43 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff1.q_ne_RNI2QSE5_LC_7_11_3 .C_ON=1'b0;
    defparam \uut.IR.ff1.q_ne_RNI2QSE5_LC_7_11_3 .SEQ_MODE=4'b0000;
    defparam \uut.IR.ff1.q_ne_RNI2QSE5_LC_7_11_3 .LUT_INIT=16'b1100100011001100;
    LogicCell40 \uut.IR.ff1.q_ne_RNI2QSE5_LC_7_11_3  (
            .in0(N__7933),
            .in1(N__5302),
            .in2(N__7975),
            .in3(N__7872),
            .lcout(\uut.ir_out_m_d_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff2.q_ne_RNI3V695_LC_7_11_4 .C_ON=1'b0;
    defparam \uut.IR.ff2.q_ne_RNI3V695_LC_7_11_4 .SEQ_MODE=4'b0000;
    defparam \uut.IR.ff2.q_ne_RNI3V695_LC_7_11_4 .LUT_INIT=16'b1111000011010000;
    LogicCell40 \uut.IR.ff2.q_ne_RNI3V695_LC_7_11_4  (
            .in0(N__7873),
            .in1(N__7934),
            .in2(N__3559),
            .in3(N__7965),
            .lcout(\uut.ir_out_m_d_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mem.data_1_0_iv_LC_7_11_6 .C_ON=1'b0;
    defparam \uut.mem.data_1_0_iv_LC_7_11_6 .SEQ_MODE=4'b0000;
    defparam \uut.mem.data_1_0_iv_LC_7_11_6 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \uut.mem.data_1_0_iv_LC_7_11_6  (
            .in0(N__6395),
            .in1(N__6349),
            .in2(N__6316),
            .in3(N__9046),
            .lcout(\uut.bus_6 ),
            .ltout(\uut.bus_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff7.q_0_ne_RNI7UKPK_LC_7_11_7 .C_ON=1'b0;
    defparam \uut.IR.ff7.q_0_ne_RNI7UKPK_LC_7_11_7 .SEQ_MODE=4'b0000;
    defparam \uut.IR.ff7.q_0_ne_RNI7UKPK_LC_7_11_7 .LUT_INIT=16'b1111001111000000;
    LogicCell40 \uut.IR.ff7.q_0_ne_RNI7UKPK_LC_7_11_7  (
            .in0(_gnd_net_),
            .in1(N__7403),
            .in2(N__3415),
            .in3(N__4042),
            .lcout(\uut.N_5_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.acc.ff5.q_RNIDGA71_LC_7_12_0 .C_ON=1'b0;
    defparam \uut.acc.ff5.q_RNIDGA71_LC_7_12_0 .SEQ_MODE=4'b0000;
    defparam \uut.acc.ff5.q_RNIDGA71_LC_7_12_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uut.acc.ff5.q_RNIDGA71_LC_7_12_0  (
            .in0(N__5878),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8271),
            .lcout(\uut.q_RNIDGA71 ),
            .ltout(\uut.q_RNIDGA71_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.b_reg.ff5.q_LC_7_12_1 .C_ON=1'b0;
    defparam \uut.b_reg.ff5.q_LC_7_12_1 .SEQ_MODE=4'b1000;
    defparam \uut.b_reg.ff5.q_LC_7_12_1 .LUT_INIT=16'b1111111111110001;
    LogicCell40 \uut.b_reg.ff5.q_LC_7_12_1  (
            .in0(N__5948),
            .in1(N__9043),
            .in2(N__3412),
            .in3(N__5905),
            .lcout(\uut.b_reg_out_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.b_reg.ff5.qC_net ),
            .ce(N__7510),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.ALU_Out_0_4_LC_7_12_2 .C_ON=1'b0;
    defparam \uut.ALU_main.ALU_Out_0_4_LC_7_12_2 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.ALU_Out_0_4_LC_7_12_2 .LUT_INIT=16'b1000100001100110;
    LogicCell40 \uut.ALU_main.ALU_Out_0_4_LC_7_12_2  (
            .in0(N__5877),
            .in1(N__3445),
            .in2(_gnd_net_),
            .in3(N__6767),
            .lcout(),
            .ltout(\uut.ALU_main.N_45_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_cry_3_c_RNIGUMDE_LC_7_12_3 .C_ON=1'b0;
    defparam \uut.ALU_main.un1_A_cry_3_c_RNIGUMDE_LC_7_12_3 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_cry_3_c_RNIGUMDE_LC_7_12_3 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \uut.ALU_main.un1_A_cry_3_c_RNIGUMDE_LC_7_12_3  (
            .in0(N__4264),
            .in1(N__6621),
            .in2(N__3409),
            .in3(N__6475),
            .lcout(\uut.alu_out_m_4 ),
            .ltout(\uut.alu_out_m_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mem.data_1_2_ivdup_LC_7_12_4 .C_ON=1'b0;
    defparam \uut.mem.data_1_2_ivdup_LC_7_12_4 .SEQ_MODE=4'b0000;
    defparam \uut.mem.data_1_2_ivdup_LC_7_12_4 .LUT_INIT=16'b1111111111110001;
    LogicCell40 \uut.mem.data_1_2_ivdup_LC_7_12_4  (
            .in0(N__9042),
            .in1(N__5947),
            .in2(N__3406),
            .in3(N__5966),
            .lcout(\uut.data_1_2_ivdup ),
            .ltout(\uut.data_1_2_ivdup_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff5.q_0_ne_RNINJRHK_LC_7_12_5 .C_ON=1'b0;
    defparam \uut.IR.ff5.q_0_ne_RNINJRHK_LC_7_12_5 .SEQ_MODE=4'b0000;
    defparam \uut.IR.ff5.q_0_ne_RNINJRHK_LC_7_12_5 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \uut.IR.ff5.q_0_ne_RNINJRHK_LC_7_12_5  (
            .in0(N__4700),
            .in1(_gnd_net_),
            .in2(N__3403),
            .in3(N__7412),
            .lcout(\uut.N_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mem.data_1_2_iv_0_LC_7_12_6 .C_ON=1'b0;
    defparam \uut.mem.data_1_2_iv_0_LC_7_12_6 .SEQ_MODE=4'b0000;
    defparam \uut.mem.data_1_2_iv_0_LC_7_12_6 .LUT_INIT=16'b1010101010101111;
    LogicCell40 \uut.mem.data_1_2_iv_0_LC_7_12_6  (
            .in0(N__5879),
            .in1(_gnd_net_),
            .in2(N__9071),
            .in3(N__5946),
            .lcout(\uut.data_1_2_iv_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_axb_4_l_ofx_LC_7_12_7 .C_ON=1'b0;
    defparam \uut.ALU_main.un1_A_axb_4_l_ofx_LC_7_12_7 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_axb_4_l_ofx_LC_7_12_7 .LUT_INIT=16'b0101010101100110;
    LogicCell40 \uut.ALU_main.un1_A_axb_4_l_ofx_LC_7_12_7  (
            .in0(N__3444),
            .in1(N__4767),
            .in2(N__5884),
            .in3(N__4419),
            .lcout(\uut.ALU_main.un1_A_axb_4_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff5.q_0_ne_LC_7_13_2 .C_ON=1'b0;
    defparam \uut.IR.ff5.q_0_ne_LC_7_13_2 .SEQ_MODE=4'b1000;
    defparam \uut.IR.ff5.q_0_ne_LC_7_13_2 .LUT_INIT=16'b1111110011111101;
    LogicCell40 \uut.IR.ff5.q_0_ne_LC_7_13_2  (
            .in0(N__5949),
            .in1(N__5906),
            .in2(N__5983),
            .in3(N__9077),
            .lcout(\uut.ir_out_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff5.q_0_neC_net ),
            .ce(N__7428),
            .sr(_gnd_net_));
    defparam \uut.seq.q_ret_RNI52E81_0_LC_7_13_3 .C_ON=1'b0;
    defparam \uut.seq.q_ret_RNI52E81_0_LC_7_13_3 .SEQ_MODE=4'b0000;
    defparam \uut.seq.q_ret_RNI52E81_0_LC_7_13_3 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uut.seq.q_ret_RNI52E81_0_LC_7_13_3  (
            .in0(N__4677),
            .in1(N__4103),
            .in2(N__3803),
            .in3(N__4022),
            .lcout(\uut.seq.q_ret_RNI52E81Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff7.q_0_ne_LC_7_13_4 .C_ON=1'b0;
    defparam \uut.IR.ff7.q_0_ne_LC_7_13_4 .SEQ_MODE=4'b1000;
    defparam \uut.IR.ff7.q_0_ne_LC_7_13_4 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \uut.IR.ff7.q_0_ne_LC_7_13_4  (
            .in0(N__6388),
            .in1(N__6359),
            .in2(N__6330),
            .in3(N__9076),
            .lcout(\uut.ir_out_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff5.q_0_neC_net ),
            .ce(N__7428),
            .sr(_gnd_net_));
    defparam \uut.IR.ff8.q_0_ne_LC_7_13_5 .C_ON=1'b0;
    defparam \uut.IR.ff8.q_0_ne_LC_7_13_5 .SEQ_MODE=4'b1000;
    defparam \uut.IR.ff8.q_0_ne_LC_7_13_5 .LUT_INIT=16'b1111110011111101;
    LogicCell40 \uut.IR.ff8.q_0_ne_LC_7_13_5  (
            .in0(N__9075),
            .in1(N__6195),
            .in2(N__6229),
            .in3(N__6885),
            .lcout(\uut.ir_out_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff5.q_0_neC_net ),
            .ce(N__7428),
            .sr(_gnd_net_));
    defparam \uut.IR.ff3.q_RNIILCK5_LC_7_14_0 .C_ON=1'b0;
    defparam \uut.IR.ff3.q_RNIILCK5_LC_7_14_0 .SEQ_MODE=4'b0000;
    defparam \uut.IR.ff3.q_RNIILCK5_LC_7_14_0 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \uut.IR.ff3.q_RNIILCK5_LC_7_14_0  (
            .in0(N__7987),
            .in1(N__7929),
            .in2(N__7254),
            .in3(N__7894),
            .lcout(),
            .ltout(\uut.ir_out_m_d_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.out_1_0_iv_2_1_LC_7_14_1 .C_ON=1'b0;
    defparam \uut.AR_BUF.out_1_0_iv_2_1_LC_7_14_1 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.out_1_0_iv_2_1_LC_7_14_1 .LUT_INIT=16'b1111111111111101;
    LogicCell40 \uut.AR_BUF.out_1_0_iv_2_1_LC_7_14_1  (
            .in0(N__3490),
            .in1(N__3436),
            .in2(N__3427),
            .in3(N__4478),
            .lcout(\uut.out_1_0_iv_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.q_ret_LC_7_14_2 .C_ON=1'b0;
    defparam \uut.seq.q_ret_LC_7_14_2 .SEQ_MODE=4'b1000;
    defparam \uut.seq.q_ret_LC_7_14_2 .LUT_INIT=16'b0000000010101010;
    LogicCell40 \uut.seq.q_ret_LC_7_14_2  (
            .in0(N__7406),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3884),
            .lcout(\uut.un1_HLT_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.seq.q_retC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.ALU_Out_0_7_LC_7_14_4 .C_ON=1'b0;
    defparam \uut.ALU_main.ALU_Out_0_7_LC_7_14_4 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.ALU_Out_0_7_LC_7_14_4 .LUT_INIT=16'b1000100001100110;
    LogicCell40 \uut.ALU_main.ALU_Out_0_7_LC_7_14_4  (
            .in0(N__4524),
            .in1(N__6177),
            .in2(_gnd_net_),
            .in3(N__6768),
            .lcout(\uut.ALU_main.N_48 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.acc.ff7.q_RNIFKC71_LC_7_14_6 .C_ON=1'b0;
    defparam \uut.acc.ff7.q_RNIFKC71_LC_7_14_6 .SEQ_MODE=4'b0000;
    defparam \uut.acc.ff7.q_RNIFKC71_LC_7_14_6 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uut.acc.ff7.q_RNIFKC71_LC_7_14_6  (
            .in0(_gnd_net_),
            .in1(N__6273),
            .in2(_gnd_net_),
            .in3(N__8272),
            .lcout(\uut.acc_out_m_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.out_1_0_iv_2_1_1_LC_7_14_7 .C_ON=1'b0;
    defparam \uut.AR_BUF.out_1_0_iv_2_1_1_LC_7_14_7 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.out_1_0_iv_2_1_1_LC_7_14_7 .LUT_INIT=16'b0011001101110111;
    LogicCell40 \uut.AR_BUF.out_1_0_iv_2_1_1_LC_7_14_7  (
            .in0(N__8375),
            .in1(N__7247),
            .in2(_gnd_net_),
            .in3(N__7139),
            .lcout(\uut.AR_BUF.out_1_0_iv_2_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff1.q_ne_LC_7_15_0 .C_ON=1'b0;
    defparam \uut.IR.ff1.q_ne_LC_7_15_0 .SEQ_MODE=4'b1000;
    defparam \uut.IR.ff1.q_ne_LC_7_15_0 .LUT_INIT=16'b1111111111110001;
    LogicCell40 \uut.IR.ff1.q_ne_LC_7_15_0  (
            .in0(N__9137),
            .in1(N__9054),
            .in2(N__9194),
            .in3(N__9239),
            .lcout(\uut.ir_out_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff1.q_neC_net ),
            .ce(N__7432),
            .sr(_gnd_net_));
    defparam \uut.IR.ff2.q_ne_LC_7_15_4 .C_ON=1'b0;
    defparam \uut.IR.ff2.q_ne_LC_7_15_4 .SEQ_MODE=4'b1000;
    defparam \uut.IR.ff2.q_ne_LC_7_15_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \uut.IR.ff2.q_ne_LC_7_15_4  (
            .in0(N__7693),
            .in1(N__7645),
            .in2(_gnd_net_),
            .in3(N__7597),
            .lcout(\uut.ir_out_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff1.q_neC_net ),
            .ce(N__7432),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_0_a5_0_2_LC_7_16_1 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_0_a5_0_2_LC_7_16_1 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_0_a5_0_2_LC_7_16_1 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \uut.AR_BUF.g0_0_a5_0_2_LC_7_16_1  (
            .in0(N__7028),
            .in1(N__7238),
            .in2(N__8716),
            .in3(N__4138),
            .lcout(),
            .ltout(\uut.AR_BUF.g0_0_a5_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_0_a5_0_LC_7_16_2 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_0_a5_0_LC_7_16_2 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_0_a5_0_LC_7_16_2 .LUT_INIT=16'b1011000010100000;
    LogicCell40 \uut.AR_BUF.g0_0_a5_0_LC_7_16_2  (
            .in0(N__4932),
            .in1(N__4702),
            .in2(N__3481),
            .in3(N__6934),
            .lcout(\uut.AR_BUF.N_9 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_1_0_1_LC_8_8_0 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_1_0_1_LC_8_8_0 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_1_0_1_LC_8_8_0 .LUT_INIT=16'b1111111110000000;
    LogicCell40 \uut.AR_BUF.g0_1_0_1_LC_8_8_0  (
            .in0(N__4044),
            .in1(N__3814),
            .in2(N__3469),
            .in3(N__3451),
            .lcout(\uut.AR_BUF.g0_1_0Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_0_o5_0_0_LC_8_8_3 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_0_o5_0_0_LC_8_8_3 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_0_o5_0_0_LC_8_8_3 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \uut.AR_BUF.g0_0_o5_0_0_LC_8_8_3  (
            .in0(N__5516),
            .in1(N__9402),
            .in2(_gnd_net_),
            .in3(N__8549),
            .lcout(\uut.AR_BUF.g0_0_o5_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_1_a10_3_0_LC_8_8_6 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_1_a10_3_0_LC_8_8_6 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_1_a10_3_0_LC_8_8_6 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uut.AR_BUF.g0_1_a10_3_0_LC_8_8_6  (
            .in0(N__5099),
            .in1(N__5357),
            .in2(N__3558),
            .in3(N__6942),
            .lcout(),
            .ltout(\uut.AR_BUF.g0_1_a10_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_1_a10_LC_8_8_7 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_1_a10_LC_8_8_7 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_1_a10_LC_8_8_7 .LUT_INIT=16'b0011000000100000;
    LogicCell40 \uut.AR_BUF.g0_1_a10_LC_8_8_7  (
            .in0(N__7032),
            .in1(N__4142),
            .in2(N__3454),
            .in3(N__4043),
            .lcout(\uut.AR_BUF.N_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_1_a10_4_LC_8_9_0 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_1_a10_4_LC_8_9_0 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_1_a10_4_LC_8_9_0 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \uut.AR_BUF.g0_1_a10_4_LC_8_9_0  (
            .in0(N__3553),
            .in1(N__4930),
            .in2(N__3943),
            .in3(N__4143),
            .lcout(),
            .ltout(\uut.AR_BUF.N_13_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_1_0_5_LC_8_9_1 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_1_0_5_LC_8_9_1 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_1_0_5_LC_8_9_1 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \uut.AR_BUF.g0_1_0_5_LC_8_9_1  (
            .in0(N__5181),
            .in1(N__3502),
            .in2(N__3604),
            .in3(N__8253),
            .lcout(),
            .ltout(\uut.AR_BUF.g0_1_0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_1_1_LC_8_9_2 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_1_1_LC_8_9_2 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_1_1_LC_8_9_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uut.AR_BUF.g0_1_1_LC_8_9_2  (
            .in0(N__3496),
            .in1(N__3565),
            .in2(N__3601),
            .in3(N__3598),
            .lcout(\uut.out_1_1_iv_3dup_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_3_a10_1_1_LC_8_9_5 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_3_a10_1_1_LC_8_9_5 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_3_a10_1_1_LC_8_9_5 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uut.AR_BUF.g0_3_a10_1_1_LC_8_9_5  (
            .in0(N__4931),
            .in1(N__8757),
            .in2(_gnd_net_),
            .in3(N__5297),
            .lcout(\uut.AR_BUF.g0_3_a10_1Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_1_0_6_LC_8_9_6 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_1_0_6_LC_8_9_6 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_1_0_6_LC_8_9_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \uut.AR_BUF.g0_1_0_6_LC_8_9_6  (
            .in0(N__3552),
            .in1(N__7760),
            .in2(N__3592),
            .in3(N__8386),
            .lcout(\uut.AR_BUF.g0_1_0_4_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_1_a8_3_LC_8_9_7 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_1_a8_3_LC_8_9_7 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_1_a8_3_LC_8_9_7 .LUT_INIT=16'b1000100000000000;
    LogicCell40 \uut.AR_BUF.g0_1_a8_3_LC_8_9_7  (
            .in0(N__9403),
            .in1(N__3551),
            .in2(_gnd_net_),
            .in3(N__8550),
            .lcout(\uut.AR_BUF.N_10 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_1_0_2_LC_8_10_0 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_1_0_2_LC_8_10_0 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_1_0_2_LC_8_10_0 .LUT_INIT=16'b1111000010000000;
    LogicCell40 \uut.AR_BUF.g0_1_0_2_LC_8_10_0  (
            .in0(N__8577),
            .in1(N__8761),
            .in2(N__5748),
            .in3(N__8657),
            .lcout(\uut.AR_BUF.g0_1_0_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.pc.program_counter_RNO_3_1_LC_8_10_1 .C_ON=1'b0;
    defparam \uut.pc.program_counter_RNO_3_1_LC_8_10_1 .SEQ_MODE=4'b0000;
    defparam \uut.pc.program_counter_RNO_3_1_LC_8_10_1 .LUT_INIT=16'b1111111111111000;
    LogicCell40 \uut.pc.program_counter_RNO_3_1_LC_8_10_1  (
            .in0(N__9401),
            .in1(N__8578),
            .in2(N__3664),
            .in3(N__7763),
            .lcout(\uut.pc.g2_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.pc.program_counter_RNO_1_1_LC_8_10_2 .C_ON=1'b0;
    defparam \uut.pc.program_counter_RNO_1_1_LC_8_10_2 .SEQ_MODE=4'b0000;
    defparam \uut.pc.program_counter_RNO_1_1_LC_8_10_2 .LUT_INIT=16'b0101101011110000;
    LogicCell40 \uut.pc.program_counter_RNO_1_1_LC_8_10_2  (
            .in0(N__5701),
            .in1(_gnd_net_),
            .in2(N__5749),
            .in3(N__7327),
            .lcout(\uut.pc.N_77_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_RNICCTC1_0_LC_8_10_3 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_RNICCTC1_0_LC_8_10_3 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_RNICCTC1_0_LC_8_10_3 .LUT_INIT=16'b1100100010001000;
    LogicCell40 \uut.seq.counter.T_1_RNICCTC1_0_LC_8_10_3  (
            .in0(N__8656),
            .in1(N__5700),
            .in2(N__8769),
            .in3(N__8576),
            .lcout(\uut.program_counter_m_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.pc.program_counter_1_LC_8_10_4 .C_ON=1'b0;
    defparam \uut.pc.program_counter_1_LC_8_10_4 .SEQ_MODE=4'b1000;
    defparam \uut.pc.program_counter_1_LC_8_10_4 .LUT_INIT=16'b1111111111100000;
    LogicCell40 \uut.pc.program_counter_1_LC_8_10_4  (
            .in0(N__7567),
            .in1(N__7643),
            .in2(N__5484),
            .in3(N__4351),
            .lcout(\uut.program_counter_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5631),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.pc.program_counter_RNO_0_0_LC_8_10_5 .C_ON=1'b0;
    defparam \uut.pc.program_counter_RNO_0_0_LC_8_10_5 .SEQ_MODE=4'b0000;
    defparam \uut.pc.program_counter_RNO_0_0_LC_8_10_5 .LUT_INIT=16'b0000000100000000;
    LogicCell40 \uut.pc.program_counter_RNO_0_0_LC_8_10_5  (
            .in0(N__9258),
            .in1(N__3610),
            .in2(N__3648),
            .in3(N__4207),
            .lcout(),
            .ltout(\uut.pc.N_4_i_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.pc.program_counter_0_LC_8_10_6 .C_ON=1'b0;
    defparam \uut.pc.program_counter_0_LC_8_10_6 .SEQ_MODE=4'b1000;
    defparam \uut.pc.program_counter_0_LC_8_10_6 .LUT_INIT=16'b0000011000000111;
    LogicCell40 \uut.pc.program_counter_0_LC_8_10_6  (
            .in0(N__5702),
            .in1(N__7328),
            .in2(N__3631),
            .in3(N__4240),
            .lcout(\uut.program_counter_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5631),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.b_reg.ff3.q_LC_8_11_1 .C_ON=1'b0;
    defparam \uut.b_reg.ff3.q_LC_8_11_1 .SEQ_MODE=4'b1000;
    defparam \uut.b_reg.ff3.q_LC_8_11_1 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \uut.b_reg.ff3.q_LC_8_11_1  (
            .in0(N__8099),
            .in1(N__3628),
            .in2(N__5451),
            .in3(N__9053),
            .lcout(\uut.b_reg_out_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.b_reg.ff3.qC_net ),
            .ce(N__7516),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.g0_1_LC_8_11_2 .C_ON=1'b0;
    defparam \uut.ALU_main.g0_1_LC_8_11_2 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.g0_1_LC_8_11_2 .LUT_INIT=16'b1000100001100110;
    LogicCell40 \uut.ALU_main.g0_1_LC_8_11_2  (
            .in0(N__4467),
            .in1(N__4499),
            .in2(_gnd_net_),
            .in3(N__6753),
            .lcout(),
            .ltout(\uut.ALU_main.N_43_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_cry_1_c_RNI46ADE_LC_8_11_3 .C_ON=1'b0;
    defparam \uut.ALU_main.un1_A_cry_1_c_RNI46ADE_LC_8_11_3 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_cry_1_c_RNI46ADE_LC_8_11_3 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \uut.ALU_main.un1_A_cry_1_c_RNI46ADE_LC_8_11_3  (
            .in0(N__6581),
            .in1(N__6463),
            .in2(N__3616),
            .in3(N__4296),
            .lcout(\uut.alu_out_m_0_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_fast_RNIVM0N3_0_LC_8_11_4 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_fast_RNIVM0N3_0_LC_8_11_4 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_fast_RNIVM0N3_0_LC_8_11_4 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uut.seq.counter.T_1_fast_RNIVM0N3_0_LC_8_11_4  (
            .in0(_gnd_net_),
            .in1(N__6752),
            .in2(_gnd_net_),
            .in3(N__4418),
            .lcout(\uut.T_1_fast_RNIVM0N3_0 ),
            .ltout(\uut.T_1_fast_RNIVM0N3_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.pc.program_counter_RNO_2_0_LC_8_11_5 .C_ON=1'b0;
    defparam \uut.pc.program_counter_RNO_2_0_LC_8_11_5 .SEQ_MODE=4'b0000;
    defparam \uut.pc.program_counter_RNO_2_0_LC_8_11_5 .LUT_INIT=16'b0101110000001100;
    LogicCell40 \uut.pc.program_counter_RNO_2_0_LC_8_11_5  (
            .in0(N__6580),
            .in1(N__4805),
            .in2(N__3613),
            .in3(N__4320),
            .lcout(\uut.pc.N_11 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_2_rep1_RNI8TE81_LC_8_12_0 .C_ON=1'b0;
    defparam \uut.seq.counter.T_2_rep1_RNI8TE81_LC_8_12_0 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_2_rep1_RNI8TE81_LC_8_12_0 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \uut.seq.counter.T_2_rep1_RNI8TE81_LC_8_12_0  (
            .in0(N__7020),
            .in1(N__4989),
            .in2(N__5100),
            .in3(N__4116),
            .lcout(),
            .ltout(\uut.seq.counter.T_2_rep1_RNI8TEZ0Z81_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_2_rep1_RNI51JC1_LC_8_12_1 .C_ON=1'b0;
    defparam \uut.seq.counter.T_2_rep1_RNI51JC1_LC_8_12_1 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_2_rep1_RNI51JC1_LC_8_12_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \uut.seq.counter.T_2_rep1_RNI51JC1_LC_8_12_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3682),
            .in3(N__3856),
            .lcout(\uut.seq.counter.un2_MAR_LD ),
            .ltout(\uut.seq.counter.un2_MAR_LD_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_RNI33MC3_3_LC_8_12_2 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_RNI33MC3_3_LC_8_12_2 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_RNI33MC3_3_LC_8_12_2 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \uut.seq.counter.T_1_RNI33MC3_3_LC_8_12_2  (
            .in0(N__5520),
            .in1(N__9395),
            .in2(N__3679),
            .in3(N__8552),
            .lcout(\uut.un1_IR_OE_4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.decoder.D_0_1_LC_8_12_3 .C_ON=1'b0;
    defparam \uut.seq.decoder.D_0_1_LC_8_12_3 .SEQ_MODE=4'b0000;
    defparam \uut.seq.decoder.D_0_1_LC_8_12_3 .LUT_INIT=16'b0101010100000000;
    LogicCell40 \uut.seq.decoder.D_0_1_LC_8_12_3  (
            .in0(N__4990),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3855),
            .lcout(\uut.D_1_0 ),
            .ltout(\uut.D_1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_RNIEDK31_2_LC_8_12_4 .C_ON=1'b0;
    defparam \uut.seq.counter.T_RNIEDK31_2_LC_8_12_4 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_RNIEDK31_2_LC_8_12_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uut.seq.counter.T_RNIEDK31_2_LC_8_12_4  (
            .in0(N__8744),
            .in1(N__4117),
            .in2(N__3676),
            .in3(N__4024),
            .lcout(\uut.un14_MAR_LD ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_2_rep1_RNI6BLF1_LC_8_12_5 .C_ON=1'b0;
    defparam \uut.seq.counter.T_2_rep1_RNI6BLF1_LC_8_12_5 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_2_rep1_RNI6BLF1_LC_8_12_5 .LUT_INIT=16'b1110111000100010;
    LogicCell40 \uut.seq.counter.T_2_rep1_RNI6BLF1_LC_8_12_5  (
            .in0(_gnd_net_),
            .in1(N__4684),
            .in2(_gnd_net_),
            .in3(N__3691),
            .lcout(\uut.T_2_rep1_RNI6BLF1 ),
            .ltout(\uut.T_2_rep1_RNI6BLF1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_RNIVVKI3_3_LC_8_12_6 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_RNIVVKI3_3_LC_8_12_6 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_RNIVVKI3_3_LC_8_12_6 .LUT_INIT=16'b0000000100000101;
    LogicCell40 \uut.seq.counter.T_1_RNIVVKI3_3_LC_8_12_6  (
            .in0(N__3673),
            .in1(N__9394),
            .in2(N__3667),
            .in3(N__8551),
            .lcout(\uut.T_1_RNIVVKI3_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.q_ret_RNI52E81_LC_8_12_7 .C_ON=1'b0;
    defparam \uut.seq.q_ret_RNI52E81_LC_8_12_7 .SEQ_MODE=4'b0000;
    defparam \uut.seq.q_ret_RNI52E81_LC_8_12_7 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \uut.seq.q_ret_RNI52E81_LC_8_12_7  (
            .in0(N__4023),
            .in1(N__3810),
            .in2(N__4136),
            .in3(N__4685),
            .lcout(\uut.un17_IR_OE_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_3_LC_8_13_0 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_3_LC_8_13_0 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_3_LC_8_13_0 .LUT_INIT=16'b1111100010001000;
    LogicCell40 \uut.AR_BUF.g0_3_LC_8_13_0  (
            .in0(N__8278),
            .in1(N__8495),
            .in2(N__8416),
            .in3(N__8359),
            .lcout(\uut.AR_BUF.g0_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff5.q_0_rep1_RNIIHI7_LC_8_13_1 .C_ON=1'b0;
    defparam \uut.IR.ff5.q_0_rep1_RNIIHI7_LC_8_13_1 .SEQ_MODE=4'b0000;
    defparam \uut.IR.ff5.q_0_rep1_RNIIHI7_LC_8_13_1 .LUT_INIT=16'b0011001111111111;
    LogicCell40 \uut.IR.ff5.q_0_rep1_RNIIHI7_LC_8_13_1  (
            .in0(_gnd_net_),
            .in1(N__5359),
            .in2(_gnd_net_),
            .in3(N__4910),
            .lcout(),
            .ltout(\uut.IR.ir_out_m_c_d_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff4.q_ne_RNINTO01_LC_8_13_2 .C_ON=1'b0;
    defparam \uut.IR.ff4.q_ne_RNINTO01_LC_8_13_2 .SEQ_MODE=4'b0000;
    defparam \uut.IR.ff4.q_ne_RNINTO01_LC_8_13_2 .LUT_INIT=16'b0000100000000000;
    LogicCell40 \uut.IR.ff4.q_ne_RNINTO01_LC_8_13_2  (
            .in0(N__8404),
            .in1(N__9460),
            .in2(N__3697),
            .in3(N__5082),
            .lcout(\uut.ir_out_m_c_d_3 ),
            .ltout(\uut.ir_out_m_c_d_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff4.q_ne_LC_8_13_3 .C_ON=1'b0;
    defparam \uut.IR.ff4.q_ne_LC_8_13_3 .SEQ_MODE=4'b1000;
    defparam \uut.IR.ff4.q_ne_LC_8_13_3 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uut.IR.ff4.q_ne_LC_8_13_3  (
            .in0(N__9808),
            .in1(N__9739),
            .in2(N__3694),
            .in3(N__9859),
            .lcout(\uut.ir_out_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff4.q_neC_net ),
            .ce(N__7401),
            .sr(_gnd_net_));
    defparam \uut.IR.ff6.q_0_ne_LC_8_13_4 .C_ON=1'b0;
    defparam \uut.IR.ff6.q_0_ne_LC_8_13_4 .SEQ_MODE=4'b1000;
    defparam \uut.IR.ff6.q_0_ne_LC_8_13_4 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \uut.IR.ff6.q_0_ne_LC_8_13_4  (
            .in0(N__6114),
            .in1(N__6141),
            .in2(N__9079),
            .in3(N__6078),
            .lcout(\uut.ir_out_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff4.q_neC_net ),
            .ce(N__7401),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_2_rep1_RNIGC8C1_LC_8_13_5 .C_ON=1'b0;
    defparam \uut.seq.counter.T_2_rep1_RNIGC8C1_LC_8_13_5 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_2_rep1_RNIGC8C1_LC_8_13_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \uut.seq.counter.T_2_rep1_RNIGC8C1_LC_8_13_5  (
            .in0(N__5081),
            .in1(N__4909),
            .in2(N__3733),
            .in3(N__4102),
            .lcout(\uut.seq.counter.T_2_rep1_RNIGC8CZ0Z1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.un13_ACC_LD_x1_LC_8_14_0 .C_ON=1'b0;
    defparam \uut.seq.un13_ACC_LD_x1_LC_8_14_0 .SEQ_MODE=4'b0000;
    defparam \uut.seq.un13_ACC_LD_x1_LC_8_14_0 .LUT_INIT=16'b0000010000000000;
    LogicCell40 \uut.seq.un13_ACC_LD_x1_LC_8_14_0  (
            .in0(N__4982),
            .in1(N__4019),
            .in2(N__4128),
            .in3(N__3849),
            .lcout(),
            .ltout(\uut.seq.un13_ACC_LD_xZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_fast_RNITEB42_0_LC_8_14_1 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_fast_RNITEB42_0_LC_8_14_1 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_fast_RNITEB42_0_LC_8_14_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \uut.seq.counter.T_1_fast_RNITEB42_0_LC_8_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__3685),
            .in3(N__4839),
            .lcout(\uut.un13_ACC_LD ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.decoder.D_6_LC_8_14_2 .C_ON=1'b0;
    defparam \uut.seq.decoder.D_6_LC_8_14_2 .SEQ_MODE=4'b0000;
    defparam \uut.seq.decoder.D_6_LC_8_14_2 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \uut.seq.decoder.D_6_LC_8_14_2  (
            .in0(N__3731),
            .in1(N__5421),
            .in2(N__5021),
            .in3(N__5349),
            .lcout(\uut.D_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff7.q_ret_1_fast_LC_8_14_3 .C_ON=1'b0;
    defparam \uut.IR.ff7.q_ret_1_fast_LC_8_14_3 .SEQ_MODE=4'b1000;
    defparam \uut.IR.ff7.q_ret_1_fast_LC_8_14_3 .LUT_INIT=16'b0101010101010101;
    LogicCell40 \uut.IR.ff7.q_ret_1_fast_LC_8_14_3  (
            .in0(N__3778),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uut.q_ret_1_fast ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff7.q_ret_1_fastC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_2_rep1_LC_8_14_4 .C_ON=1'b0;
    defparam \uut.seq.counter.T_2_rep1_LC_8_14_4 .SEQ_MODE=4'b1000;
    defparam \uut.seq.counter.T_2_rep1_LC_8_14_4 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uut.seq.counter.T_2_rep1_LC_8_14_4  (
            .in0(N__7405),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uut.T_2_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff7.q_ret_1_fastC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.q_ret_RNIAFH51_LC_8_14_5 .C_ON=1'b0;
    defparam \uut.seq.q_ret_RNIAFH51_LC_8_14_5 .SEQ_MODE=4'b0000;
    defparam \uut.seq.q_ret_RNIAFH51_LC_8_14_5 .LUT_INIT=16'b0000000010000000;
    LogicCell40 \uut.seq.q_ret_RNIAFH51_LC_8_14_5  (
            .in0(N__4020),
            .in1(N__3797),
            .in2(N__5358),
            .in3(N__4101),
            .lcout(\uut.un17_IR_OE ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff7.q_ret_1_LC_8_14_6 .C_ON=1'b0;
    defparam \uut.IR.ff7.q_ret_1_LC_8_14_6 .SEQ_MODE=4'b1000;
    defparam \uut.IR.ff7.q_ret_1_LC_8_14_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uut.IR.ff7.q_ret_1_LC_8_14_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3777),
            .lcout(\uut.ir_out_i_2_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff7.q_ret_1_fastC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff7.q_0_fast_LC_8_14_7 .C_ON=1'b0;
    defparam \uut.IR.ff7.q_0_fast_LC_8_14_7 .SEQ_MODE=4'b1000;
    defparam \uut.IR.ff7.q_0_fast_LC_8_14_7 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uut.IR.ff7.q_0_fast_LC_8_14_7  (
            .in0(N__4021),
            .in1(N__3760),
            .in2(_gnd_net_),
            .in3(N__7404),
            .lcout(\uut.q_0_fast ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff7.q_ret_1_fastC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff5.q_0_rep1_LC_8_15_0 .C_ON=1'b0;
    defparam \uut.IR.ff5.q_0_rep1_LC_8_15_0 .SEQ_MODE=4'b1000;
    defparam \uut.IR.ff5.q_0_rep1_LC_8_15_0 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uut.IR.ff5.q_0_rep1_LC_8_15_0  (
            .in0(N__7419),
            .in1(N__3709),
            .in2(_gnd_net_),
            .in3(N__4704),
            .lcout(\uut.ir_out_4_rep1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff5.q_0_rep1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff8.q_0_fast_LC_8_15_1 .C_ON=1'b0;
    defparam \uut.IR.ff8.q_0_fast_LC_8_15_1 .SEQ_MODE=4'b1000;
    defparam \uut.IR.ff8.q_0_fast_LC_8_15_1 .LUT_INIT=16'b1011101110001000;
    LogicCell40 \uut.IR.ff8.q_0_fast_LC_8_15_1  (
            .in0(N__3748),
            .in1(N__7420),
            .in2(_gnd_net_),
            .in3(N__4135),
            .lcout(\uut.q_0_fast_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff5.q_0_rep1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.decoder.D_2_0_x_LC_8_15_2 .C_ON=1'b0;
    defparam \uut.seq.decoder.D_2_0_x_LC_8_15_2 .SEQ_MODE=4'b0000;
    defparam \uut.seq.decoder.D_2_0_x_LC_8_15_2 .LUT_INIT=16'b0001000100000000;
    LogicCell40 \uut.seq.decoder.D_2_0_x_LC_8_15_2  (
            .in0(N__4978),
            .in1(N__5419),
            .in2(_gnd_net_),
            .in3(N__4869),
            .lcout(),
            .ltout(\uut.seq.D_2_0_x_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_fast_RNI874E2_0_LC_8_15_3 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_fast_RNI874E2_0_LC_8_15_3 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_fast_RNI874E2_0_LC_8_15_3 .LUT_INIT=16'b1110110000000000;
    LogicCell40 \uut.seq.counter.T_1_fast_RNI874E2_0_LC_8_15_3  (
            .in0(N__5012),
            .in1(N__4782),
            .in2(N__3736),
            .in3(N__4841),
            .lcout(\uut.S0_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff6.q_ret_1_fast_LC_8_15_4 .C_ON=1'b0;
    defparam \uut.IR.ff6.q_ret_1_fast_LC_8_15_4 .SEQ_MODE=4'b1000;
    defparam \uut.IR.ff6.q_ret_1_fast_LC_8_15_4 .LUT_INIT=16'b0011001100110011;
    LogicCell40 \uut.IR.ff6.q_ret_1_fast_LC_8_15_4  (
            .in0(_gnd_net_),
            .in1(N__3891),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uut.q_ret_1_fast_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff5.q_0_rep1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.decoder.D_4_0_LC_8_15_5 .C_ON=1'b0;
    defparam \uut.seq.decoder.D_4_0_LC_8_15_5 .SEQ_MODE=4'b0000;
    defparam \uut.seq.decoder.D_4_0_LC_8_15_5 .LUT_INIT=16'b0001000000000000;
    LogicCell40 \uut.seq.decoder.D_4_0_LC_8_15_5  (
            .in0(N__5420),
            .in1(N__4977),
            .in2(N__3732),
            .in3(N__3848),
            .lcout(\uut.seq.D_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff5.q_0_fast_LC_8_15_6 .C_ON=1'b0;
    defparam \uut.IR.ff5.q_0_fast_LC_8_15_6 .SEQ_MODE=4'b1000;
    defparam \uut.IR.ff5.q_0_fast_LC_8_15_6 .LUT_INIT=16'b1101110110001000;
    LogicCell40 \uut.IR.ff5.q_0_fast_LC_8_15_6  (
            .in0(N__7418),
            .in1(N__3708),
            .in2(_gnd_net_),
            .in3(N__4703),
            .lcout(\uut.ir_out_fast_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff5.q_0_rep1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_2_LC_8_15_7 .C_ON=1'b0;
    defparam \uut.seq.counter.T_2_LC_8_15_7 .SEQ_MODE=4'b1000;
    defparam \uut.seq.counter.T_2_LC_8_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut.seq.counter.T_2_LC_8_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7421),
            .lcout(\uut.T_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff5.q_0_rep1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_fast_3_LC_8_16_0 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_fast_3_LC_8_16_0 .SEQ_MODE=4'b1000;
    defparam \uut.seq.counter.T_1_fast_3_LC_8_16_0 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uut.seq.counter.T_1_fast_3_LC_8_16_0  (
            .in0(N__8715),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uut.seq.counter.T_1_fastZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.seq.counter.T_1_fast_3C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_fast_RNI4JTR1_0_LC_8_16_1 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_fast_RNI4JTR1_0_LC_8_16_1 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_fast_RNI4JTR1_0_LC_8_16_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uut.seq.counter.T_1_fast_RNI4JTR1_0_LC_8_16_1  (
            .in0(N__7029),
            .in1(N__6935),
            .in2(N__7059),
            .in3(N__4843),
            .lcout(),
            .ltout(\uut.seq.counter.un4_ACC_LD_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_RNI4F1C2_3_LC_8_16_2 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_RNI4F1C2_3_LC_8_16_2 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_RNI4F1C2_3_LC_8_16_2 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \uut.seq.counter.T_1_RNI4F1C2_3_LC_8_16_2  (
            .in0(N__9469),
            .in1(N__3979),
            .in2(N__3910),
            .in3(N__9396),
            .lcout(\uut.seq.counter.ACC_LD_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff6.q_ret_1_LC_8_16_6 .C_ON=1'b0;
    defparam \uut.IR.ff6.q_ret_1_LC_8_16_6 .SEQ_MODE=4'b1000;
    defparam \uut.IR.ff6.q_ret_1_LC_8_16_6 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uut.IR.ff6.q_ret_1_LC_8_16_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__3892),
            .lcout(\uut.ir_out_i_2_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.seq.counter.T_1_fast_3C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_fast_RNI6J9S_3_LC_8_16_7 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_fast_RNI6J9S_3_LC_8_16_7 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_fast_RNI6J9S_3_LC_8_16_7 .LUT_INIT=16'b0000000011110111;
    LogicCell40 \uut.seq.counter.T_1_fast_RNI6J9S_3_LC_8_16_7  (
            .in0(N__4641),
            .in1(N__3847),
            .in2(N__4988),
            .in3(N__9419),
            .lcout(\uut.seq.counter.T_1_fast_RNI6J9SZ0Z_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_3_3_LC_9_8_1 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_3_3_LC_9_8_1 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_3_3_LC_9_8_1 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \uut.AR_BUF.g0_3_3_LC_9_8_1  (
            .in0(N__4201),
            .in1(N__3958),
            .in2(N__5245),
            .in3(N__8286),
            .lcout(\uut.AR_BUF.g0_3Z0Z_3 ),
            .ltout(\uut.AR_BUF.g0_3Z0Z_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.acc.ff1.q_LC_9_8_2 .C_ON=1'b0;
    defparam \uut.acc.ff1.q_LC_9_8_2 .SEQ_MODE=4'b1000;
    defparam \uut.acc.ff1.q_LC_9_8_2 .LUT_INIT=16'b1111101011111011;
    LogicCell40 \uut.acc.ff1.q_LC_9_8_2  (
            .in0(N__9220),
            .in1(N__9139),
            .in2(N__3826),
            .in3(N__9078),
            .lcout(\uut.acc_out_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.acc.ff1.qC_net ),
            .ce(N__5841),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.out_1_2_iv_1_LC_9_8_4 .C_ON=1'b0;
    defparam \uut.AR_BUF.out_1_2_iv_1_LC_9_8_4 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.out_1_2_iv_1_LC_9_8_4 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \uut.AR_BUF.out_1_2_iv_1_LC_9_8_4  (
            .in0(N__3949),
            .in1(N__5237),
            .in2(_gnd_net_),
            .in3(N__4200),
            .lcout(\uut.AR_BUF.out_1_2_ivZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_3_a10_0_2_LC_9_9_1 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_3_a10_0_2_LC_9_9_1 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_3_a10_0_2_LC_9_9_1 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uut.AR_BUF.g0_3_a10_0_2_LC_9_9_1  (
            .in0(N__5300),
            .in1(N__4144),
            .in2(N__8773),
            .in3(N__4045),
            .lcout(),
            .ltout(\uut.AR_BUF.g0_3_a10_0Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_3_0_LC_9_9_2 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_3_0_LC_9_9_2 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_3_0_LC_9_9_2 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \uut.AR_BUF.g0_3_0_LC_9_9_2  (
            .in0(N__3985),
            .in1(N__3978),
            .in2(N__3961),
            .in3(N__9468),
            .lcout(\uut.AR_BUF.g0_3Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff1.q_ne_RNIKEQ11_LC_9_9_4 .C_ON=1'b0;
    defparam \uut.IR.ff1.q_ne_RNIKEQ11_LC_9_9_4 .SEQ_MODE=4'b0000;
    defparam \uut.IR.ff1.q_ne_RNIKEQ11_LC_9_9_4 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uut.IR.ff1.q_ne_RNIKEQ11_LC_9_9_4  (
            .in0(_gnd_net_),
            .in1(N__5301),
            .in2(_gnd_net_),
            .in3(N__7140),
            .lcout(),
            .ltout(\uut.ir_out_m_c_d_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.out_1_2_iv_2_LC_9_9_5 .C_ON=1'b0;
    defparam \uut.AR_BUF.out_1_2_iv_2_LC_9_9_5 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.out_1_2_iv_2_LC_9_9_5 .LUT_INIT=16'b1111111011111100;
    LogicCell40 \uut.AR_BUF.out_1_2_iv_2_LC_9_9_5  (
            .in0(N__3925),
            .in1(N__4225),
            .in2(N__3952),
            .in3(N__7761),
            .lcout(\uut.AR_BUF.out_1_2_ivZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_1_a10_4_1_LC_9_9_7 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_1_a10_4_1_LC_9_9_7 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_1_a10_4_1_LC_9_9_7 .LUT_INIT=16'b1100110000000000;
    LogicCell40 \uut.AR_BUF.g0_1_a10_4_1_LC_9_9_7  (
            .in0(_gnd_net_),
            .in1(N__5101),
            .in2(_gnd_net_),
            .in3(N__7033),
            .lcout(\uut.AR_BUF.g0_1_a10_4Z0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_3_2_LC_9_10_0 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_3_2_LC_9_10_0 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_3_2_LC_9_10_0 .LUT_INIT=16'b1111111110001000;
    LogicCell40 \uut.AR_BUF.g0_3_2_LC_9_10_0  (
            .in0(N__7759),
            .in1(N__3924),
            .in2(_gnd_net_),
            .in3(N__4224),
            .lcout(),
            .ltout(\uut.AR_BUF.g0_3Z0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_3_6_LC_9_10_1 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_3_6_LC_9_10_1 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_3_6_LC_9_10_1 .LUT_INIT=16'b1111110011111110;
    LogicCell40 \uut.AR_BUF.g0_3_6_LC_9_10_1  (
            .in0(N__5299),
            .in1(N__4183),
            .in2(N__3931),
            .in3(N__7893),
            .lcout(\uut.AR_BUF.g0_3Z0Z_6 ),
            .ltout(\uut.AR_BUF.g0_3Z0Z_6_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR.ff1.q_ne_LC_9_10_2 .C_ON=1'b0;
    defparam \uut.AR.ff1.q_ne_LC_9_10_2 .SEQ_MODE=4'b1000;
    defparam \uut.AR.ff1.q_ne_LC_9_10_2 .LUT_INIT=16'b1111101011111011;
    LogicCell40 \uut.AR.ff1.q_ne_LC_9_10_2  (
            .in0(N__9175),
            .in1(N__9138),
            .in2(N__3928),
            .in3(N__9037),
            .lcout(\uut.AR_out_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.AR.ff1.q_neC_net ),
            .ce(N__8027),
            .sr(_gnd_net_));
    defparam \uut.pc.program_counter_RNO_3_0_LC_9_10_3 .C_ON=1'b0;
    defparam \uut.pc.program_counter_RNO_3_0_LC_9_10_3 .SEQ_MODE=4'b0000;
    defparam \uut.pc.program_counter_RNO_3_0_LC_9_10_3 .LUT_INIT=16'b1111100011111111;
    LogicCell40 \uut.pc.program_counter_RNO_3_0_LC_9_10_3  (
            .in0(N__3923),
            .in1(N__7758),
            .in2(N__7360),
            .in3(N__5206),
            .lcout(),
            .ltout(\uut.pc.G_26_i_a4_5_sx_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.pc.program_counter_RNO_1_0_LC_9_10_4 .C_ON=1'b0;
    defparam \uut.pc.program_counter_RNO_1_0_LC_9_10_4 .SEQ_MODE=4'b0000;
    defparam \uut.pc.program_counter_RNO_1_0_LC_9_10_4 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uut.pc.program_counter_RNO_1_0_LC_9_10_4  (
            .in0(N__4239),
            .in1(N__4223),
            .in2(N__4210),
            .in3(N__4194),
            .lcout(\uut.pc.G_26_i_a4_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff1.q_ne_RNIMP2B1_LC_9_10_5 .C_ON=1'b0;
    defparam \uut.IR.ff1.q_ne_RNIMP2B1_LC_9_10_5 .SEQ_MODE=4'b0000;
    defparam \uut.IR.ff1.q_ne_RNIMP2B1_LC_9_10_5 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uut.IR.ff1.q_ne_RNIMP2B1_LC_9_10_5  (
            .in0(N__5298),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8360),
            .lcout(\uut.ir_out_m_c_c_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_fast_RNIFJ9BG_0_LC_9_10_6 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_fast_RNIFJ9BG_0_LC_9_10_6 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_fast_RNIFJ9BG_0_LC_9_10_6 .LUT_INIT=16'b0010111000100010;
    LogicCell40 \uut.seq.counter.T_1_fast_RNIFJ9BG_0_LC_9_10_6  (
            .in0(N__4806),
            .in1(N__6467),
            .in2(N__6603),
            .in3(N__4326),
            .lcout(\uut.alu_out_m_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_fast_RNIFJ9BG_0_0_LC_9_10_7 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_fast_RNIFJ9BG_0_0_LC_9_10_7 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_fast_RNIFJ9BG_0_0_LC_9_10_7 .LUT_INIT=16'b0000101011001100;
    LogicCell40 \uut.seq.counter.T_1_fast_RNIFJ9BG_0_0_LC_9_10_7  (
            .in0(N__4327),
            .in1(N__4807),
            .in2(N__6610),
            .in3(N__6474),
            .lcout(\uut.alu_out_m_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_axb_3_l_ofx_LC_9_11_0 .C_ON=1'b0;
    defparam \uut.ALU_main.un1_A_axb_3_l_ofx_LC_9_11_0 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_axb_3_l_ofx_LC_9_11_0 .LUT_INIT=16'b0011001101100110;
    LogicCell40 \uut.ALU_main.un1_A_axb_3_l_ofx_LC_9_11_0  (
            .in0(N__4760),
            .in1(N__6653),
            .in2(N__8497),
            .in3(N__4416),
            .lcout(\uut.ALU_main.un1_A_axb_3_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.b_reg.ff4.q_LC_9_11_1 .C_ON=1'b0;
    defparam \uut.b_reg.ff4.q_LC_9_11_1 .SEQ_MODE=4'b1000;
    defparam \uut.b_reg.ff4.q_LC_9_11_1 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uut.b_reg.ff4.q_LC_9_11_1  (
            .in0(N__9850),
            .in1(N__9802),
            .in2(N__9771),
            .in3(N__9713),
            .lcout(\uut.b_reg_out_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.b_reg.ff4.qC_net ),
            .ce(N__7487),
            .sr(_gnd_net_));
    defparam \uut.pc.program_counter_RNO_4_1_LC_9_11_4 .C_ON=1'b0;
    defparam \uut.pc.program_counter_RNO_4_1_LC_9_11_4 .SEQ_MODE=4'b0000;
    defparam \uut.pc.program_counter_RNO_4_1_LC_9_11_4 .LUT_INIT=16'b1001001010000000;
    LogicCell40 \uut.pc.program_counter_RNO_4_1_LC_9_11_4  (
            .in0(N__7549),
            .in1(N__6754),
            .in2(N__5192),
            .in3(N__4417),
            .lcout(),
            .ltout(\uut.pc.program_counter_4_a1_0_0_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.pc.program_counter_RNO_2_1_LC_9_11_5 .C_ON=1'b0;
    defparam \uut.pc.program_counter_RNO_2_1_LC_9_11_5 .SEQ_MODE=4'b0000;
    defparam \uut.pc.program_counter_RNO_2_1_LC_9_11_5 .LUT_INIT=16'b1111010011110000;
    LogicCell40 \uut.pc.program_counter_RNO_2_1_LC_9_11_5  (
            .in0(N__6582),
            .in1(N__6456),
            .in2(N__4162),
            .in3(N__5124),
            .lcout(),
            .ltout(\uut.pc.g1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.pc.program_counter_RNO_0_1_LC_9_11_6 .C_ON=1'b0;
    defparam \uut.pc.program_counter_RNO_0_1_LC_9_11_6 .SEQ_MODE=4'b0000;
    defparam \uut.pc.program_counter_RNO_0_1_LC_9_11_6 .LUT_INIT=16'b1100110011100100;
    LogicCell40 \uut.pc.program_counter_RNO_0_1_LC_9_11_6  (
            .in0(N__4159),
            .in1(N__4153),
            .in2(N__4147),
            .in3(N__7386),
            .lcout(\uut.pc.program_counter_0_1_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_fast_RNI6RIE3_0_LC_9_11_7 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_fast_RNI6RIE3_0_LC_9_11_7 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_fast_RNI6RIE3_0_LC_9_11_7 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uut.seq.counter.T_1_fast_RNI6RIE3_0_LC_9_11_7  (
            .in0(_gnd_net_),
            .in1(N__4627),
            .in2(_gnd_net_),
            .in3(N__4759),
            .lcout(\uut.un1_ALU_en_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_cry_0_c_THRU_CRY_0_LC_9_12_0 .C_ON=1'b1;
    defparam \uut.ALU_main.un1_A_cry_0_c_THRU_CRY_0_LC_9_12_0 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_cry_0_c_THRU_CRY_0_LC_9_12_0 .LUT_INIT=16'b0000000000000000;
    LogicCell40 \uut.ALU_main.un1_A_cry_0_c_THRU_CRY_0_LC_9_12_0  (
            .in0(_gnd_net_),
            .in1(N__4341),
            .in2(N__4345),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_9_12_0_),
            .carryout(\uut.ALU_main.un1_A_cry_0_c_THRU_CO ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_cry_0_s_LC_9_12_1 .C_ON=1'b1;
    defparam \uut.ALU_main.un1_A_cry_0_s_LC_9_12_1 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_cry_0_s_LC_9_12_1 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uut.ALU_main.un1_A_cry_0_s_LC_9_12_1  (
            .in0(_gnd_net_),
            .in1(N__5243),
            .in2(N__4534),
            .in3(N__4309),
            .lcout(\uut.un1_A_cry_0_s ),
            .ltout(),
            .carryin(\uut.ALU_main.un1_A_cry_0_c_THRU_CO ),
            .carryout(\uut.ALU_main.un1_A_cry_0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_cry_0_c_RNI3CH45_LC_9_12_2 .C_ON=1'b1;
    defparam \uut.ALU_main.un1_A_cry_0_c_RNI3CH45_LC_9_12_2 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_cry_0_c_RNI3CH45_LC_9_12_2 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uut.ALU_main.un1_A_cry_0_c_RNI3CH45_LC_9_12_2  (
            .in0(_gnd_net_),
            .in1(N__4588),
            .in2(N__5193),
            .in3(N__4306),
            .lcout(\uut.un1_A_cry_0_c_RNI3CH45 ),
            .ltout(),
            .carryin(\uut.ALU_main.un1_A_cry_0 ),
            .carryout(\uut.ALU_main.un1_A_cry_1 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_cry_1_c_RNI7KL45_LC_9_12_3 .C_ON=1'b1;
    defparam \uut.ALU_main.un1_A_cry_1_c_RNI7KL45_LC_9_12_3 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_cry_1_c_RNI7KL45_LC_9_12_3 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uut.ALU_main.un1_A_cry_1_c_RNI7KL45_LC_9_12_3  (
            .in0(_gnd_net_),
            .in1(N__4357),
            .in2(N__4479),
            .in3(N__4285),
            .lcout(\uut.ALU_main.un1_A_cry_1_c_RNI7KLZ0Z45 ),
            .ltout(),
            .carryin(\uut.ALU_main.un1_A_cry_1 ),
            .carryout(\uut.ALU_main.un1_A_cry_2_cZ0 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_cry_2_c_RNIBSP45_LC_9_12_4 .C_ON=1'b1;
    defparam \uut.ALU_main.un1_A_cry_2_c_RNIBSP45_LC_9_12_4 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_cry_2_c_RNIBSP45_LC_9_12_4 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uut.ALU_main.un1_A_cry_2_c_RNIBSP45_LC_9_12_4  (
            .in0(_gnd_net_),
            .in1(N__4282),
            .in2(N__8496),
            .in3(N__4276),
            .lcout(\uut.un1_A_cry_2_c_RNIBSP45 ),
            .ltout(),
            .carryin(\uut.ALU_main.un1_A_cry_2_cZ0 ),
            .carryout(\uut.ALU_main.un1_A_cry_3 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_cry_3_c_RNIF4U45_LC_9_12_5 .C_ON=1'b1;
    defparam \uut.ALU_main.un1_A_cry_3_c_RNIF4U45_LC_9_12_5 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_cry_3_c_RNIF4U45_LC_9_12_5 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uut.ALU_main.un1_A_cry_3_c_RNIF4U45_LC_9_12_5  (
            .in0(_gnd_net_),
            .in1(N__4273),
            .in2(N__5883),
            .in3(N__4255),
            .lcout(\uut.ALU_main.un1_A_cry_3_c_RNIF4UZ0Z45 ),
            .ltout(),
            .carryin(\uut.ALU_main.un1_A_cry_3 ),
            .carryout(\uut.ALU_main.un1_A_cry_4 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_cry_4_c_RNIJC255_LC_9_12_6 .C_ON=1'b1;
    defparam \uut.ALU_main.un1_A_cry_4_c_RNIJC255_LC_9_12_6 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_cry_4_c_RNIJC255_LC_9_12_6 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uut.ALU_main.un1_A_cry_4_c_RNIJC255_LC_9_12_6  (
            .in0(_gnd_net_),
            .in1(N__4540),
            .in2(N__6028),
            .in3(N__4243),
            .lcout(\uut.ALU_main.un1_A_cry_4_c_RNIJCZ0Z255 ),
            .ltout(),
            .carryin(\uut.ALU_main.un1_A_cry_4 ),
            .carryout(\uut.ALU_main.un1_A_cry_5 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_cry_5_c_RNINK655_LC_9_12_7 .C_ON=1'b1;
    defparam \uut.ALU_main.un1_A_cry_5_c_RNINK655_LC_9_12_7 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_cry_5_c_RNINK655_LC_9_12_7 .LUT_INIT=16'b1100001100111100;
    LogicCell40 \uut.ALU_main.un1_A_cry_5_c_RNINK655_LC_9_12_7  (
            .in0(_gnd_net_),
            .in1(N__4564),
            .in2(N__6274),
            .in3(N__4603),
            .lcout(\uut.ALU_main.un1_A_cry_5_c_RNINKZ0Z655 ),
            .ltout(),
            .carryin(\uut.ALU_main.un1_A_cry_5 ),
            .carryout(\uut.ALU_main.un1_A_cry_6 ),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_cry_6_c_RNINIMN4_LC_9_13_0 .C_ON=1'b0;
    defparam \uut.ALU_main.un1_A_cry_6_c_RNINIMN4_LC_9_13_0 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_cry_6_c_RNINIMN4_LC_9_13_0 .LUT_INIT=16'b0011001111001100;
    LogicCell40 \uut.ALU_main.un1_A_cry_6_c_RNINIMN4_LC_9_13_0  (
            .in0(_gnd_net_),
            .in1(N__4510),
            .in2(_gnd_net_),
            .in3(N__4600),
            .lcout(\uut.ALU_main.un1_A_cry_6_c_RNINIMNZ0Z4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_axb_1_l_ofx_LC_9_13_1 .C_ON=1'b0;
    defparam \uut.ALU_main.un1_A_axb_1_l_ofx_LC_9_13_1 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_axb_1_l_ofx_LC_9_13_1 .LUT_INIT=16'b0101010101100110;
    LogicCell40 \uut.ALU_main.un1_A_axb_1_l_ofx_LC_9_13_1  (
            .in0(N__7548),
            .in1(N__4737),
            .in2(N__5194),
            .in3(N__4396),
            .lcout(\uut.ALU_main.un1_A_axb_1_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_axb_6_l_ofx_LC_9_13_2 .C_ON=1'b0;
    defparam \uut.ALU_main.un1_A_axb_6_l_ofx_LC_9_13_2 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_axb_6_l_ofx_LC_9_13_2 .LUT_INIT=16'b0000010111111010;
    LogicCell40 \uut.ALU_main.un1_A_axb_6_l_ofx_LC_9_13_2  (
            .in0(N__4399),
            .in1(N__6265),
            .in2(N__4757),
            .in3(N__4581),
            .lcout(\uut.ALU_main.un1_A_axb_6_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_axb_5_l_ofx_LC_9_13_3 .C_ON=1'b0;
    defparam \uut.ALU_main.un1_A_axb_5_l_ofx_LC_9_13_3 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_axb_5_l_ofx_LC_9_13_3 .LUT_INIT=16'b0101010101100110;
    LogicCell40 \uut.ALU_main.un1_A_axb_5_l_ofx_LC_9_13_3  (
            .in0(N__4558),
            .in1(N__4739),
            .in2(N__6031),
            .in3(N__4398),
            .lcout(\uut.ALU_main.un1_A_axb_5_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_axb_0_l_ofx_LC_9_13_5 .C_ON=1'b0;
    defparam \uut.ALU_main.un1_A_axb_0_l_ofx_LC_9_13_5 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_axb_0_l_ofx_LC_9_13_5 .LUT_INIT=16'b0011001100111100;
    LogicCell40 \uut.ALU_main.un1_A_axb_0_l_ofx_LC_9_13_5  (
            .in0(N__5244),
            .in1(N__6798),
            .in2(N__4415),
            .in3(N__4736),
            .lcout(\uut.ALU_main.un1_A_axb_0_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_axb_7_LC_9_13_6 .C_ON=1'b0;
    defparam \uut.ALU_main.un1_A_axb_7_LC_9_13_6 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_axb_7_LC_9_13_6 .LUT_INIT=16'b1100100100110110;
    LogicCell40 \uut.ALU_main.un1_A_axb_7_LC_9_13_6  (
            .in0(N__4400),
            .in1(N__4525),
            .in2(N__4758),
            .in3(N__6170),
            .lcout(\uut.ALU_main.un1_A_axbZ0Z_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_axb_2_l_ofx_LC_9_13_7 .C_ON=1'b0;
    defparam \uut.ALU_main.un1_A_axb_2_l_ofx_LC_9_13_7 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_axb_2_l_ofx_LC_9_13_7 .LUT_INIT=16'b0101010101100110;
    LogicCell40 \uut.ALU_main.un1_A_axb_2_l_ofx_LC_9_13_7  (
            .in0(N__4504),
            .in1(N__4738),
            .in2(N__4480),
            .in3(N__4397),
            .lcout(\uut.ALU_main.un1_A_axb_2_l_ofxZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_2_rep1_RNIJDGJ_LC_9_14_0 .C_ON=1'b0;
    defparam \uut.seq.counter.T_2_rep1_RNIJDGJ_LC_9_14_0 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_2_rep1_RNIJDGJ_LC_9_14_0 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uut.seq.counter.T_2_rep1_RNIJDGJ_LC_9_14_0  (
            .in0(N__5414),
            .in1(N__5339),
            .in2(N__5092),
            .in3(N__4906),
            .lcout(),
            .ltout(\uut.seq.counter.T_2_rep1_RNIJDGJZ0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_2_rep1_RNIHU2O_LC_9_14_1 .C_ON=1'b0;
    defparam \uut.seq.counter.T_2_rep1_RNIHU2O_LC_9_14_1 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_2_rep1_RNIHU2O_LC_9_14_1 .LUT_INIT=16'b1111000010101010;
    LogicCell40 \uut.seq.counter.T_2_rep1_RNIHU2O_LC_9_14_1  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__4786),
            .in3(N__4865),
            .lcout(\uut.un11_MAR_LD ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.B_LD_2_tz_LC_9_14_2 .C_ON=1'b0;
    defparam \uut.seq.B_LD_2_tz_LC_9_14_2 .SEQ_MODE=4'b0000;
    defparam \uut.seq.B_LD_2_tz_LC_9_14_2 .LUT_INIT=16'b0001001100110011;
    LogicCell40 \uut.seq.B_LD_2_tz_LC_9_14_2  (
            .in0(N__9458),
            .in1(N__4783),
            .in2(N__5029),
            .in3(N__5341),
            .lcout(\uut.B_LD_0_2_tz ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.decoder.D_0_2_LC_9_14_3 .C_ON=1'b0;
    defparam \uut.seq.decoder.D_0_2_LC_9_14_3 .SEQ_MODE=4'b0000;
    defparam \uut.seq.decoder.D_0_2_LC_9_14_3 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \uut.seq.decoder.D_0_2_LC_9_14_3  (
            .in0(_gnd_net_),
            .in1(N__4863),
            .in2(_gnd_net_),
            .in3(N__5413),
            .lcout(\uut.D_1_3 ),
            .ltout(\uut.D_1_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_fast_RNI28LI1_0_0_LC_9_14_4 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_fast_RNI28LI1_0_0_LC_9_14_4 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_fast_RNI28LI1_0_0_LC_9_14_4 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uut.seq.counter.T_1_fast_RNI28LI1_0_0_LC_9_14_4  (
            .in0(N__4840),
            .in1(N__5340),
            .in2(N__4771),
            .in3(N__4907),
            .lcout(\uut.un7_ACC_LD ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_2_rep1_RNIJ9B11_LC_9_14_5 .C_ON=1'b0;
    defparam \uut.seq.counter.T_2_rep1_RNIJ9B11_LC_9_14_5 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_2_rep1_RNIJ9B11_LC_9_14_5 .LUT_INIT=16'b1100110010101010;
    LogicCell40 \uut.seq.counter.T_2_rep1_RNIJ9B11_LC_9_14_5  (
            .in0(N__5047),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__5415),
            .lcout(\uut.un5_MAR_LD ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.decoder.D_2_0_LC_9_14_6 .C_ON=1'b0;
    defparam \uut.seq.decoder.D_2_0_LC_9_14_6 .SEQ_MODE=4'b0000;
    defparam \uut.seq.decoder.D_2_0_LC_9_14_6 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \uut.seq.decoder.D_2_0_LC_9_14_6  (
            .in0(N__4864),
            .in1(N__4981),
            .in2(N__5028),
            .in3(N__5422),
            .lcout(\uut.seq.D_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_RNIEPQK_2_LC_9_14_7 .C_ON=1'b0;
    defparam \uut.seq.counter.T_RNIEPQK_2_LC_9_14_7 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_RNIEPQK_2_LC_9_14_7 .LUT_INIT=16'b0010000000000000;
    LogicCell40 \uut.seq.counter.T_RNIEPQK_2_LC_9_14_7  (
            .in0(N__4908),
            .in1(N__4705),
            .in2(N__8717),
            .in3(N__9459),
            .lcout(\uut.un8_MAR_LD ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_fast_RNIU5S31_0_LC_9_15_1 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_fast_RNIU5S31_0_LC_9_15_1 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_fast_RNIU5S31_0_LC_9_15_1 .LUT_INIT=16'b0000000000000001;
    LogicCell40 \uut.seq.counter.T_1_fast_RNIU5S31_0_LC_9_15_1  (
            .in0(N__9420),
            .in1(N__4642),
            .in2(N__5377),
            .in3(N__4996),
            .lcout(\uut.seq.counter.T_4 ),
            .ltout(\uut.seq.counter.T_4_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_fast_RNI4JTR1_0_0_LC_9_15_2 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_fast_RNI4JTR1_0_0_LC_9_15_2 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_fast_RNI4JTR1_0_0_LC_9_15_2 .LUT_INIT=16'b0111111111111111;
    LogicCell40 \uut.seq.counter.T_1_fast_RNI4JTR1_0_0_LC_9_15_2  (
            .in0(N__7049),
            .in1(N__7019),
            .in2(N__4630),
            .in3(N__6927),
            .lcout(\uut.seq.counter.T_1_fast_RNI4JTR1_0Z0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_2_rep1_RNIV9NU_LC_9_15_3 .C_ON=1'b0;
    defparam \uut.seq.counter.T_2_rep1_RNIV9NU_LC_9_15_3 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_2_rep1_RNIV9NU_LC_9_15_3 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uut.seq.counter.T_2_rep1_RNIV9NU_LC_9_15_3  (
            .in0(N__6926),
            .in1(N__5080),
            .in2(N__7031),
            .in3(N__4980),
            .lcout(\uut.seq.counter.T_2_rep1_RNIV9NUZ0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.IR.ff6.q_0_fast_LC_9_15_4 .C_ON=1'b0;
    defparam \uut.IR.ff6.q_0_fast_LC_9_15_4 .SEQ_MODE=4'b1000;
    defparam \uut.IR.ff6.q_0_fast_LC_9_15_4 .LUT_INIT=16'b1010101011001100;
    LogicCell40 \uut.IR.ff6.q_0_fast_LC_9_15_4  (
            .in0(N__5041),
            .in1(N__4929),
            .in2(_gnd_net_),
            .in3(N__7416),
            .lcout(\uut.q_0_fast_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff6.q_0_fastC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_fast_2_LC_9_15_5 .C_ON=1'b0;
    defparam \uut.seq.counter.T_fast_2_LC_9_15_5 .SEQ_MODE=4'b1000;
    defparam \uut.seq.counter.T_fast_2_LC_9_15_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uut.seq.counter.T_fast_2_LC_9_15_5  (
            .in0(N__7417),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uut.seq.counter.T_fastZ0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff6.q_0_fastC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_fast_1_LC_9_15_6 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_fast_1_LC_9_15_6 .SEQ_MODE=4'b1000;
    defparam \uut.seq.counter.T_1_fast_1_LC_9_15_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut.seq.counter.T_1_fast_1_LC_9_15_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8658),
            .lcout(\uut.seq.counter.T_1_fastZ0Z_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff6.q_0_fastC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_fast_0_LC_9_15_7 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_fast_0_LC_9_15_7 .SEQ_MODE=4'b1000;
    defparam \uut.seq.counter.T_1_fast_0_LC_9_15_7 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut.seq.counter.T_1_fast_0_LC_9_15_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7837),
            .lcout(\uut.seq.counter.T_1_fastZ0Z_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff6.q_0_fastC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.decoder.D_1_0_2_LC_9_16_0 .C_ON=1'b0;
    defparam \uut.seq.decoder.D_1_0_2_LC_9_16_0 .SEQ_MODE=4'b0000;
    defparam \uut.seq.decoder.D_1_0_2_LC_9_16_0 .LUT_INIT=16'b0000000011001100;
    LogicCell40 \uut.seq.decoder.D_1_0_2_LC_9_16_0  (
            .in0(_gnd_net_),
            .in1(N__4979),
            .in2(_gnd_net_),
            .in3(N__5417),
            .lcout(\uut.seq.D_2_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.un10_ACC_LD_x1_LC_9_16_1 .C_ON=1'b0;
    defparam \uut.seq.un10_ACC_LD_x1_LC_9_16_1 .SEQ_MODE=4'b0000;
    defparam \uut.seq.un10_ACC_LD_x1_LC_9_16_1 .LUT_INIT=16'b0100000000000000;
    LogicCell40 \uut.seq.un10_ACC_LD_x1_LC_9_16_1  (
            .in0(N__5418),
            .in1(N__4928),
            .in2(N__5356),
            .in3(N__4870),
            .lcout(),
            .ltout(\uut.seq.un10_ACC_LD_xZ0Z1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_fast_RNI28LI1_0_LC_9_16_2 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_fast_RNI28LI1_0_LC_9_16_2 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_fast_RNI28LI1_0_LC_9_16_2 .LUT_INIT=16'b1110001011100010;
    LogicCell40 \uut.seq.counter.T_1_fast_RNI28LI1_0_LC_9_16_2  (
            .in0(_gnd_net_),
            .in1(N__4842),
            .in2(N__4813),
            .in3(_gnd_net_),
            .lcout(\uut.T_1_fast_RNI28LI1_0 ),
            .ltout(\uut.T_1_fast_RNI28LI1_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.ALU_Out_0_0_LC_9_16_3 .C_ON=1'b0;
    defparam \uut.ALU_main.ALU_Out_0_0_LC_9_16_3 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.ALU_Out_0_0_LC_9_16_3 .LUT_INIT=16'b1010010100001010;
    LogicCell40 \uut.ALU_main.ALU_Out_0_0_LC_9_16_3  (
            .in0(N__5242),
            .in1(_gnd_net_),
            .in2(N__4810),
            .in3(N__6799),
            .lcout(\uut.N_41 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_fast_RNIH09P_2_LC_9_16_4 .C_ON=1'b0;
    defparam \uut.seq.counter.T_fast_RNIH09P_2_LC_9_16_4 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_fast_RNIH09P_2_LC_9_16_4 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uut.seq.counter.T_fast_RNIH09P_2_LC_9_16_4  (
            .in0(N__6925),
            .in1(N__5416),
            .in2(N__7030),
            .in3(N__5376),
            .lcout(),
            .ltout(\uut.seq.counter.T_fast_RNIH09PZ0Z_2_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_fast_RNICCPP_2_LC_9_16_5 .C_ON=1'b0;
    defparam \uut.seq.counter.T_fast_RNICCPP_2_LC_9_16_5 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_fast_RNICCPP_2_LC_9_16_5 .LUT_INIT=16'b1010101011110000;
    LogicCell40 \uut.seq.counter.T_fast_RNICCPP_2_LC_9_16_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__5362),
            .in3(N__5342),
            .lcout(\uut.OUT_LD ),
            .ltout(\uut.OUT_LD_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.pc.program_counter_RNO_4_0_LC_9_16_6 .C_ON=1'b0;
    defparam \uut.pc.program_counter_RNO_4_0_LC_9_16_6 .SEQ_MODE=4'b0000;
    defparam \uut.pc.program_counter_RNO_4_0_LC_9_16_6 .LUT_INIT=16'b0001010100111111;
    LogicCell40 \uut.pc.program_counter_RNO_4_0_LC_9_16_6  (
            .in0(N__5283),
            .in1(N__5241),
            .in2(N__5209),
            .in3(N__7132),
            .lcout(\uut.pc.G_26_i_a4_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.ALU_Out_0_1_LC_11_9_0 .C_ON=1'b0;
    defparam \uut.ALU_main.ALU_Out_0_1_LC_11_9_0 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.ALU_Out_0_1_LC_11_9_0 .LUT_INIT=16'b1001100101000100;
    LogicCell40 \uut.ALU_main.ALU_Out_0_1_LC_11_9_0  (
            .in0(N__6773),
            .in1(N__5182),
            .in2(_gnd_net_),
            .in3(N__7547),
            .lcout(),
            .ltout(\uut.ALU_main.ALU_Out_0Z0Z_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_cry_0_c_RNIUP3DE_LC_11_9_1 .C_ON=1'b0;
    defparam \uut.ALU_main.un1_A_cry_0_c_RNIUP3DE_LC_11_9_1 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_cry_0_c_RNIUP3DE_LC_11_9_1 .LUT_INIT=16'b0111010000110000;
    LogicCell40 \uut.ALU_main.un1_A_cry_0_c_RNIUP3DE_LC_11_9_1  (
            .in0(N__6617),
            .in1(N__6500),
            .in2(N__5134),
            .in3(N__5131),
            .lcout(\uut.alu_out_m_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_4_LC_11_9_6 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_4_LC_11_9_6 .SEQ_MODE=4'b1000;
    defparam \uut.seq.counter.T_1_4_LC_11_9_6 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut.seq.counter.T_1_4_LC_11_9_6  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__9393),
            .lcout(\uut.seq.counter.T_1Z0Z_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.seq.counter.T_1_4C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.g0_0_LC_11_9_7 .C_ON=1'b0;
    defparam \uut.ALU_main.g0_0_LC_11_9_7 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.g0_0_LC_11_9_7 .LUT_INIT=16'b1000100001100110;
    LogicCell40 \uut.ALU_main.g0_0_LC_11_9_7  (
            .in0(N__8488),
            .in1(N__6672),
            .in2(_gnd_net_),
            .in3(N__6772),
            .lcout(\uut.ALU_main.N_44_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_RNI215E1_0_LC_11_10_0 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_RNI215E1_0_LC_11_10_0 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_RNI215E1_0_LC_11_10_0 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uut.seq.counter.T_1_RNI215E1_0_LC_11_10_0  (
            .in0(_gnd_net_),
            .in1(N__5113),
            .in2(_gnd_net_),
            .in3(N__8654),
            .lcout(\uut.seq.counter.MAR_LD_0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.pc.program_counter_RNO_3_3_LC_11_10_1 .C_ON=1'b0;
    defparam \uut.pc.program_counter_RNO_3_3_LC_11_10_1 .SEQ_MODE=4'b0000;
    defparam \uut.pc.program_counter_RNO_3_3_LC_11_10_1 .LUT_INIT=16'b1000000000000000;
    LogicCell40 \uut.pc.program_counter_RNO_3_3_LC_11_10_1  (
            .in0(N__5793),
            .in1(N__7308),
            .in2(N__5763),
            .in3(N__5709),
            .lcout(\uut.pc.g1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.pc.g0_2_LC_11_10_2 .C_ON=1'b0;
    defparam \uut.pc.g0_2_LC_11_10_2 .SEQ_MODE=4'b0000;
    defparam \uut.pc.g0_2_LC_11_10_2 .LUT_INIT=16'b0101010100010001;
    LogicCell40 \uut.pc.g0_2_LC_11_10_2  (
            .in0(N__7309),
            .in1(N__5494),
            .in2(_gnd_net_),
            .in3(N__7779),
            .lcout(\uut.pc.un1_inc_0_0 ),
            .ltout(\uut.pc.un1_inc_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.pc.program_counter_RNO_1_3_LC_11_10_3 .C_ON=1'b0;
    defparam \uut.pc.program_counter_RNO_1_3_LC_11_10_3 .SEQ_MODE=4'b0000;
    defparam \uut.pc.program_counter_RNO_1_3_LC_11_10_3 .LUT_INIT=16'b1111001111111100;
    LogicCell40 \uut.pc.program_counter_RNO_1_3_LC_11_10_3  (
            .in0(_gnd_net_),
            .in1(N__5530),
            .in2(N__5524),
            .in3(N__8602),
            .lcout(\uut.pc.g0_rn_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_1_LC_11_10_4 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_1_LC_11_10_4 .SEQ_MODE=4'b1000;
    defparam \uut.seq.counter.T_1_1_LC_11_10_4 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut.seq.counter.T_1_1_LC_11_10_4  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8655),
            .lcout(\uut.inc ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.seq.counter.T_1_1C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_RNIU1302_3_LC_11_10_5 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_RNIU1302_3_LC_11_10_5 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_RNIU1302_3_LC_11_10_5 .LUT_INIT=16'b0001000100110011;
    LogicCell40 \uut.seq.counter.T_1_RNIU1302_3_LC_11_10_5  (
            .in0(N__9400),
            .in1(N__5521),
            .in2(_gnd_net_),
            .in3(N__8574),
            .lcout(\uut.PC_LD_0_0 ),
            .ltout(\uut.PC_LD_0_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.pc.un1_inc_LC_11_10_6 .C_ON=1'b0;
    defparam \uut.pc.un1_inc_LC_11_10_6 .SEQ_MODE=4'b0000;
    defparam \uut.pc.un1_inc_LC_11_10_6 .LUT_INIT=16'b0101010100000101;
    LogicCell40 \uut.pc.un1_inc_LC_11_10_6  (
            .in0(N__7310),
            .in1(_gnd_net_),
            .in2(N__5488),
            .in3(N__7780),
            .lcout(\uut.pc.un1_inc_0 ),
            .ltout(\uut.pc.un1_inc_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.pc.program_counter_RNO_0_2_LC_11_10_7 .C_ON=1'b0;
    defparam \uut.pc.program_counter_RNO_0_2_LC_11_10_7 .SEQ_MODE=4'b0000;
    defparam \uut.pc.program_counter_RNO_0_2_LC_11_10_7 .LUT_INIT=16'b0000001101010011;
    LogicCell40 \uut.pc.program_counter_RNO_0_2_LC_11_10_7  (
            .in0(N__7209),
            .in1(N__5680),
            .in2(N__5464),
            .in3(N__9032),
            .lcout(\uut.pc.program_counter_4_1_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mem.data_2_7_0__m13_LC_11_11_0 .C_ON=1'b0;
    defparam \uut.mem.data_2_7_0__m13_LC_11_11_0 .SEQ_MODE=4'b0000;
    defparam \uut.mem.data_2_7_0__m13_LC_11_11_0 .LUT_INIT=16'b0111111110011011;
    LogicCell40 \uut.mem.data_2_7_0__m13_LC_11_11_0  (
            .in0(N__8851),
            .in1(N__9607),
            .in2(N__9676),
            .in3(N__9525),
            .lcout(\uut.m13 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mar.ff2.q_ne_LC_11_11_1 .C_ON=1'b0;
    defparam \uut.mar.ff2.q_ne_LC_11_11_1 .SEQ_MODE=4'b1000;
    defparam \uut.mar.ff2.q_ne_LC_11_11_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \uut.mar.ff2.q_ne_LC_11_11_1  (
            .in0(N__7680),
            .in1(N__7636),
            .in2(_gnd_net_),
            .in3(N__7589),
            .lcout(\uut.mar_out_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.mar.ff2.q_neC_net ),
            .ce(N__8799),
            .sr(_gnd_net_));
    defparam \uut.mem.data_2_7_0__m20_LC_11_11_2 .C_ON=1'b0;
    defparam \uut.mem.data_2_7_0__m20_LC_11_11_2 .SEQ_MODE=4'b0000;
    defparam \uut.mem.data_2_7_0__m20_LC_11_11_2 .LUT_INIT=16'b0011110111011111;
    LogicCell40 \uut.mem.data_2_7_0__m20_LC_11_11_2  (
            .in0(N__8848),
            .in1(N__9600),
            .in2(N__9675),
            .in3(N__9522),
            .lcout(\uut.mem.m20 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mem.data_2_7_0__m22_LC_11_11_3 .C_ON=1'b0;
    defparam \uut.mem.data_2_7_0__m22_LC_11_11_3 .SEQ_MODE=4'b0000;
    defparam \uut.mem.data_2_7_0__m22_LC_11_11_3 .LUT_INIT=16'b0111001101110111;
    LogicCell40 \uut.mem.data_2_7_0__m22_LC_11_11_3  (
            .in0(N__9524),
            .in1(N__9670),
            .in2(N__9613),
            .in3(N__8850),
            .lcout(\uut.mem.N_29_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mem.data_2_7_0__m18_LC_11_11_5 .C_ON=1'b0;
    defparam \uut.mem.data_2_7_0__m18_LC_11_11_5 .SEQ_MODE=4'b0000;
    defparam \uut.mem.data_2_7_0__m18_LC_11_11_5 .LUT_INIT=16'b0111011101100101;
    LogicCell40 \uut.mem.data_2_7_0__m18_LC_11_11_5  (
            .in0(N__9523),
            .in1(N__9671),
            .in2(N__9612),
            .in3(N__8849),
            .lcout(\uut.mem.i2_mux ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.pc.program_counter_RNO_1_2_LC_11_11_7 .C_ON=1'b0;
    defparam \uut.pc.program_counter_RNO_1_2_LC_11_11_7 .SEQ_MODE=4'b0000;
    defparam \uut.pc.program_counter_RNO_1_2_LC_11_11_7 .LUT_INIT=16'b0110101010101010;
    LogicCell40 \uut.pc.program_counter_RNO_1_2_LC_11_11_7  (
            .in0(N__5797),
            .in1(N__7311),
            .in2(N__5767),
            .in3(N__5713),
            .lcout(\uut.pc.program_counter_RNO_1Z0Z_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mem.data_2_7_0__g0_0_LC_11_12_0 .C_ON=1'b0;
    defparam \uut.mem.data_2_7_0__g0_0_LC_11_12_0 .SEQ_MODE=4'b0000;
    defparam \uut.mem.data_2_7_0__g0_0_LC_11_12_0 .LUT_INIT=16'b0110101111101111;
    LogicCell40 \uut.mem.data_2_7_0__g0_0_LC_11_12_0  (
            .in0(N__9520),
            .in1(N__8846),
            .in2(N__9610),
            .in3(N__9654),
            .lcout(\uut.N_14_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.g0_LC_11_12_1 .C_ON=1'b0;
    defparam \uut.ALU_main.g0_LC_11_12_1 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.g0_LC_11_12_1 .LUT_INIT=16'b1000100001100110;
    LogicCell40 \uut.ALU_main.g0_LC_11_12_1  (
            .in0(N__8464),
            .in1(N__6668),
            .in2(_gnd_net_),
            .in3(N__6761),
            .lcout(),
            .ltout(\uut.N_44_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.pc.program_counter_RNO_0_3_LC_11_12_2 .C_ON=1'b0;
    defparam \uut.pc.program_counter_RNO_0_3_LC_11_12_2 .SEQ_MODE=4'b0000;
    defparam \uut.pc.program_counter_RNO_0_3_LC_11_12_2 .LUT_INIT=16'b0111001001010000;
    LogicCell40 \uut.pc.program_counter_RNO_0_3_LC_11_12_2  (
            .in0(N__6497),
            .in1(N__6622),
            .in2(N__5674),
            .in3(N__6635),
            .lcout(),
            .ltout(\uut.pc.alu_out_m_0_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.pc.program_counter_3_LC_11_12_3 .C_ON=1'b0;
    defparam \uut.pc.program_counter_3_LC_11_12_3 .SEQ_MODE=4'b1000;
    defparam \uut.pc.program_counter_3_LC_11_12_3 .LUT_INIT=16'b1111110010101010;
    LogicCell40 \uut.pc.program_counter_3_LC_11_12_3  (
            .in0(N__5671),
            .in1(N__7810),
            .in2(N__5662),
            .in3(N__7843),
            .lcout(\uut.program_counter_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__5648),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mem.data_2_7_0__g0_LC_11_12_4 .C_ON=1'b0;
    defparam \uut.mem.data_2_7_0__g0_LC_11_12_4 .SEQ_MODE=4'b0000;
    defparam \uut.mem.data_2_7_0__g0_LC_11_12_4 .LUT_INIT=16'b0010101010100000;
    LogicCell40 \uut.mem.data_2_7_0__g0_LC_11_12_4  (
            .in0(N__9521),
            .in1(N__8847),
            .in2(N__9611),
            .in3(N__9655),
            .lcout(\uut.N_16_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_cry_2_c_RNIAIGDE_LC_11_12_5 .C_ON=1'b0;
    defparam \uut.ALU_main.un1_A_cry_2_c_RNIAIGDE_LC_11_12_5 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_cry_2_c_RNIAIGDE_LC_11_12_5 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \uut.ALU_main.un1_A_cry_2_c_RNIAIGDE_LC_11_12_5  (
            .in0(N__6636),
            .in1(N__6614),
            .in2(N__5542),
            .in3(N__6498),
            .lcout(\uut.alu_out_m_1_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.ALU_Out_0_3_LC_11_12_6 .C_ON=1'b0;
    defparam \uut.ALU_main.ALU_Out_0_3_LC_11_12_6 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.ALU_Out_0_3_LC_11_12_6 .LUT_INIT=16'b1010010101010000;
    LogicCell40 \uut.ALU_main.ALU_Out_0_3_LC_11_12_6  (
            .in0(N__6762),
            .in1(_gnd_net_),
            .in2(N__6673),
            .in3(N__8465),
            .lcout(),
            .ltout(\uut.ALU_main.N_44_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.ALU_main.un1_A_cry_2_c_RNIAIGDE_0_LC_11_12_7 .C_ON=1'b0;
    defparam \uut.ALU_main.un1_A_cry_2_c_RNIAIGDE_0_LC_11_12_7 .SEQ_MODE=4'b0000;
    defparam \uut.ALU_main.un1_A_cry_2_c_RNIAIGDE_0_LC_11_12_7 .LUT_INIT=16'b0010001011110000;
    LogicCell40 \uut.ALU_main.un1_A_cry_2_c_RNIAIGDE_0_LC_11_12_7  (
            .in0(N__6637),
            .in1(N__6615),
            .in2(N__6505),
            .in3(N__6499),
            .lcout(\uut.alu_out_m_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.acc.ff4.q_LC_11_13_0 .C_ON=1'b0;
    defparam \uut.acc.ff4.q_LC_11_13_0 .SEQ_MODE=4'b1000;
    defparam \uut.acc.ff4.q_LC_11_13_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uut.acc.ff4.q_LC_11_13_0  (
            .in0(N__9804),
            .in1(N__9852),
            .in2(N__9763),
            .in3(N__9718),
            .lcout(\uut.acc_out_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.acc.ff4.qC_net ),
            .ce(N__5837),
            .sr(_gnd_net_));
    defparam \uut.acc.ff7.q_LC_11_13_1 .C_ON=1'b0;
    defparam \uut.acc.ff7.q_LC_11_13_1 .SEQ_MODE=4'b1000;
    defparam \uut.acc.ff7.q_LC_11_13_1 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \uut.acc.ff7.q_LC_11_13_1  (
            .in0(N__6406),
            .in1(N__6367),
            .in2(N__6320),
            .in3(N__8975),
            .lcout(\uut.acc_out_6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.acc.ff4.qC_net ),
            .ce(N__5837),
            .sr(_gnd_net_));
    defparam \uut.acc.ff8.q_LC_11_13_2 .C_ON=1'b0;
    defparam \uut.acc.ff8.q_LC_11_13_2 .SEQ_MODE=4'b1000;
    defparam \uut.acc.ff8.q_LC_11_13_2 .LUT_INIT=16'b1111111111001101;
    LogicCell40 \uut.acc.ff8.q_LC_11_13_2  (
            .in0(N__8972),
            .in1(N__6228),
            .in2(N__6884),
            .in3(N__6199),
            .lcout(\uut.acc_out_7 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.acc.ff4.qC_net ),
            .ce(N__5837),
            .sr(_gnd_net_));
    defparam \uut.acc.ff6.q_LC_11_13_3 .C_ON=1'b0;
    defparam \uut.acc.ff6.q_LC_11_13_3 .SEQ_MODE=4'b1000;
    defparam \uut.acc.ff6.q_LC_11_13_3 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \uut.acc.ff6.q_LC_11_13_3  (
            .in0(N__6145),
            .in1(N__6115),
            .in2(N__6070),
            .in3(N__8974),
            .lcout(\uut.acc_out_5 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.acc.ff4.qC_net ),
            .ce(N__5837),
            .sr(_gnd_net_));
    defparam \uut.acc.ff5.q_LC_11_13_4 .C_ON=1'b0;
    defparam \uut.acc.ff5.q_LC_11_13_4 .SEQ_MODE=4'b1000;
    defparam \uut.acc.ff5.q_LC_11_13_4 .LUT_INIT=16'b1111111111001101;
    LogicCell40 \uut.acc.ff5.q_LC_11_13_4  (
            .in0(N__8973),
            .in1(N__5979),
            .in2(N__5953),
            .in3(N__5917),
            .lcout(\uut.acc_out_4 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.acc.ff4.qC_net ),
            .ce(N__5837),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_RNIFRTJ2_3_LC_11_14_0 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_RNIFRTJ2_3_LC_11_14_0 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_RNIFRTJ2_3_LC_11_14_0 .LUT_INIT=16'b0100010011001100;
    LogicCell40 \uut.seq.counter.T_1_RNIFRTJ2_3_LC_11_14_0  (
            .in0(N__9279),
            .in1(N__9363),
            .in2(_gnd_net_),
            .in3(N__9310),
            .lcout(\uut.B_LD_0_i ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.B_LD_1_tz_LC_11_14_1 .C_ON=1'b0;
    defparam \uut.seq.B_LD_1_tz_LC_11_14_1 .SEQ_MODE=4'b0000;
    defparam \uut.seq.B_LD_1_tz_LC_11_14_1 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \uut.seq.B_LD_1_tz_LC_11_14_1  (
            .in0(N__7060),
            .in1(N__7027),
            .in2(N__6955),
            .in3(N__6943),
            .lcout(\uut.B_LD_0_1_tz ),
            .ltout(\uut.B_LD_0_1_tz_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_RNII3T14_3_LC_11_14_2 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_RNII3T14_3_LC_11_14_2 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_RNII3T14_3_LC_11_14_2 .LUT_INIT=16'b1011001100000000;
    LogicCell40 \uut.seq.counter.T_1_RNII3T14_3_LC_11_14_2  (
            .in0(N__9278),
            .in1(N__9362),
            .in2(N__6892),
            .in3(N__9297),
            .lcout(\uut.ROM_OE ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mem.data_2_7_0__m26_LC_11_14_3 .C_ON=1'b0;
    defparam \uut.mem.data_2_7_0__m26_LC_11_14_3 .SEQ_MODE=4'b0000;
    defparam \uut.mem.data_2_7_0__m26_LC_11_14_3 .LUT_INIT=16'b0111011001101101;
    LogicCell40 \uut.mem.data_2_7_0__m26_LC_11_14_3  (
            .in0(N__8843),
            .in1(N__9589),
            .in2(N__9544),
            .in3(N__9653),
            .lcout(\uut.mem.i2_mux_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.out_reg.ff3.q_LC_11_14_4 .C_ON=1'b0;
    defparam \uut.out_reg.ff3.q_LC_11_14_4 .SEQ_MODE=4'b1000;
    defparam \uut.out_reg.ff3.q_LC_11_14_4 .LUT_INIT=16'b1110111011110000;
    LogicCell40 \uut.out_reg.ff3.q_LC_11_14_4  (
            .in0(N__8077),
            .in1(N__6847),
            .in2(N__6834),
            .in3(N__8280),
            .lcout(LED3_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.out_reg.ff3.qC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_3_LC_11_14_5 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_3_LC_11_14_5 .SEQ_MODE=4'b1000;
    defparam \uut.seq.counter.T_1_3_LC_11_14_5 .LUT_INIT=16'b1010101010101010;
    LogicCell40 \uut.seq.counter.T_1_3_LC_11_14_5  (
            .in0(N__8768),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(\uut.T_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.out_reg.ff3.qC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mem.data_2_7_0__m10_LC_11_14_6 .C_ON=1'b0;
    defparam \uut.mem.data_2_7_0__m10_LC_11_14_6 .SEQ_MODE=4'b0000;
    defparam \uut.mem.data_2_7_0__m10_LC_11_14_6 .LUT_INIT=16'b0111101111001111;
    LogicCell40 \uut.mem.data_2_7_0__m10_LC_11_14_6  (
            .in0(N__9652),
            .in1(N__9539),
            .in2(N__9608),
            .in3(N__8842),
            .lcout(\uut.m10 ),
            .ltout(\uut.m10_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mem.data_2_7_0__N_11_i_m_LC_11_14_7 .C_ON=1'b0;
    defparam \uut.mem.data_2_7_0__N_11_i_m_LC_11_14_7 .SEQ_MODE=4'b0000;
    defparam \uut.mem.data_2_7_0__N_11_i_m_LC_11_14_7 .LUT_INIT=16'b0000000000001111;
    LogicCell40 \uut.mem.data_2_7_0__N_11_i_m_LC_11_14_7  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__6802),
            .in3(N__8923),
            .lcout(\uut.N_11_i_m ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.b_reg.ff1.q_LC_11_15_0 .C_ON=1'b0;
    defparam \uut.b_reg.ff1.q_LC_11_15_0 .SEQ_MODE=4'b1000;
    defparam \uut.b_reg.ff1.q_LC_11_15_0 .LUT_INIT=16'b1111101011111011;
    LogicCell40 \uut.b_reg.ff1.q_LC_11_15_0  (
            .in0(N__9240),
            .in1(N__9123),
            .in2(N__9195),
            .in3(N__8976),
            .lcout(\uut.b_reg_out_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.b_reg.ff1.qC_net ),
            .ce(N__7481),
            .sr(_gnd_net_));
    defparam \uut.b_reg.ff2.q_LC_11_15_1 .C_ON=1'b0;
    defparam \uut.b_reg.ff2.q_LC_11_15_1 .SEQ_MODE=4'b1000;
    defparam \uut.b_reg.ff2.q_LC_11_15_1 .LUT_INIT=16'b1111111111101110;
    LogicCell40 \uut.b_reg.ff2.q_LC_11_15_1  (
            .in0(N__7688),
            .in1(N__7623),
            .in2(_gnd_net_),
            .in3(N__7596),
            .lcout(\uut.b_reg_out_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.b_reg.ff1.qC_net ),
            .ce(N__7481),
            .sr(_gnd_net_));
    defparam \uut.IR.ff3.q_LC_11_16_0 .C_ON=1'b0;
    defparam \uut.IR.ff3.q_LC_11_16_0 .SEQ_MODE=4'b1000;
    defparam \uut.IR.ff3.q_LC_11_16_0 .LUT_INIT=16'b1111101011001100;
    LogicCell40 \uut.IR.ff3.q_LC_11_16_0  (
            .in0(N__8073),
            .in1(N__7237),
            .in2(N__8125),
            .in3(N__7402),
            .lcout(\uut.ir_out_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.IR.ff3.qC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_RNI3K4S_2_LC_12_10_0 .C_ON=1'b0;
    defparam \uut.seq.counter.T_RNI3K4S_2_LC_12_10_0 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_RNI3K4S_2_LC_12_10_0 .LUT_INIT=16'b1010101000000000;
    LogicCell40 \uut.seq.counter.T_RNI3K4S_2_LC_12_10_0  (
            .in0(N__8575),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8767),
            .lcout(\uut.AR_LD ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_9_LC_12_10_2 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_9_LC_12_10_2 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_9_LC_12_10_2 .LUT_INIT=16'b1111111100010001;
    LogicCell40 \uut.AR_BUF.g0_9_LC_12_10_2  (
            .in0(N__7210),
            .in1(N__9033),
            .in2(_gnd_net_),
            .in3(N__7192),
            .lcout(\uut.out_1_0_iv_3 ),
            .ltout(\uut.out_1_0_iv_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR.ff3.q_LC_12_10_3 .C_ON=1'b0;
    defparam \uut.AR.ff3.q_LC_12_10_3 .SEQ_MODE=4'b1000;
    defparam \uut.AR.ff3.q_LC_12_10_3 .LUT_INIT=16'b1111110110101000;
    LogicCell40 \uut.AR.ff3.q_LC_12_10_3  (
            .in0(N__8023),
            .in1(N__8108),
            .in2(N__7174),
            .in3(N__7163),
            .lcout(\uut.AR_out_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.AR.ff3.qC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_2_rep1_RNI48EP1_LC_12_10_6 .C_ON=1'b0;
    defparam \uut.seq.counter.T_2_rep1_RNI48EP1_LC_12_10_6 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_2_rep1_RNI48EP1_LC_12_10_6 .LUT_INIT=16'b0000000000110011;
    LogicCell40 \uut.seq.counter.T_2_rep1_RNI48EP1_LC_12_10_6  (
            .in0(_gnd_net_),
            .in1(N__8384),
            .in2(_gnd_net_),
            .in3(N__7141),
            .lcout(\uut.MAR_LD_1 ),
            .ltout(\uut.MAR_LD_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_RNI2G205_0_LC_12_10_7 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_RNI2G205_0_LC_12_10_7 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_RNI2G205_0_LC_12_10_7 .LUT_INIT=16'b0000000000100000;
    LogicCell40 \uut.seq.counter.T_1_RNI2G205_0_LC_12_10_7  (
            .in0(N__7090),
            .in1(N__7986),
            .in2(N__7084),
            .in3(N__7939),
            .lcout(\uut.MAR_LD_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_5_LC_12_11_1 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_5_LC_12_11_1 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_5_LC_12_11_1 .LUT_INIT=16'b1111111111001101;
    LogicCell40 \uut.AR_BUF.g0_5_LC_12_11_1  (
            .in0(N__8985),
            .in1(N__7699),
            .in2(N__7081),
            .in3(N__7072),
            .lcout(\uut.AR_BUF.g0Z0Z_5 ),
            .ltout(\uut.AR_BUF.g0Z0Z_5_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR.ff4.q_ne_LC_12_11_2 .C_ON=1'b0;
    defparam \uut.AR.ff4.q_ne_LC_12_11_2 .SEQ_MODE=4'b1000;
    defparam \uut.AR.ff4.q_ne_LC_12_11_2 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uut.AR.ff4.q_ne_LC_12_11_2  (
            .in0(N__9712),
            .in1(N__9767),
            .in2(N__7063),
            .in3(N__9836),
            .lcout(\uut.AR_out_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.AR.ff4.q_neC_net ),
            .ce(N__8031),
            .sr(_gnd_net_));
    defparam \uut.IR.ff4.q_ne_RNI59RD5_LC_12_11_3 .C_ON=1'b0;
    defparam \uut.IR.ff4.q_ne_RNI59RD5_LC_12_11_3 .SEQ_MODE=4'b0000;
    defparam \uut.IR.ff4.q_ne_RNI59RD5_LC_12_11_3 .LUT_INIT=16'b1110000011110000;
    LogicCell40 \uut.IR.ff4.q_ne_RNI59RD5_LC_12_11_3  (
            .in0(N__7985),
            .in1(N__7935),
            .in2(N__8431),
            .in3(N__7892),
            .lcout(\uut.ir_out_m_d_3 ),
            .ltout(\uut.ir_out_m_d_3_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.pc.program_counter_RNO_2_3_LC_12_11_4 .C_ON=1'b0;
    defparam \uut.pc.program_counter_RNO_2_3_LC_12_11_4 .SEQ_MODE=4'b0000;
    defparam \uut.pc.program_counter_RNO_2_3_LC_12_11_4 .LUT_INIT=16'b0000000000001100;
    LogicCell40 \uut.pc.program_counter_RNO_2_3_LC_12_11_4  (
            .in0(_gnd_net_),
            .in1(N__7852),
            .in2(N__7846),
            .in3(N__8301),
            .lcout(\uut.pc.g0_sn ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.out_1_iv_2_LC_12_11_5 .C_ON=1'b0;
    defparam \uut.AR_BUF.out_1_iv_2_LC_12_11_5 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.out_1_iv_2_LC_12_11_5 .LUT_INIT=16'b1111111011101110;
    LogicCell40 \uut.AR_BUF.out_1_iv_2_LC_12_11_5  (
            .in0(N__8503),
            .in1(N__9711),
            .in2(N__7803),
            .in3(N__7781),
            .lcout(\uut.out_1_iv_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_0_LC_12_12_2 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_0_LC_12_12_2 .SEQ_MODE=4'b1000;
    defparam \uut.seq.counter.T_1_0_LC_12_12_2 .LUT_INIT=16'b1111111100000000;
    LogicCell40 \uut.seq.counter.T_1_0_LC_12_12_2  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__7836),
            .lcout(\uut.T_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.seq.counter.T_1_0C_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.out_1_ivdup_0_LC_12_12_3 .C_ON=1'b0;
    defparam \uut.AR_BUF.out_1_ivdup_0_LC_12_12_3 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.out_1_ivdup_0_LC_12_12_3 .LUT_INIT=16'b1110110010100000;
    LogicCell40 \uut.AR_BUF.out_1_ivdup_0_LC_12_12_3  (
            .in0(N__8261),
            .in1(N__8426),
            .in2(N__8478),
            .in3(N__8383),
            .lcout(),
            .ltout(\uut.AR_BUF.out_1_ivdupZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_0_LC_12_12_4 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_0_LC_12_12_4 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_0_LC_12_12_4 .LUT_INIT=16'b1111000011110111;
    LogicCell40 \uut.AR_BUF.g0_0_LC_12_12_4  (
            .in0(N__9865),
            .in1(N__9526),
            .in2(N__7813),
            .in3(N__8984),
            .lcout(\uut.g0_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_RNI0KMT_0_LC_12_12_5 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_RNI0KMT_0_LC_12_12_5 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_RNI0KMT_0_LC_12_12_5 .LUT_INIT=16'b1110111011001100;
    LogicCell40 \uut.seq.counter.T_1_RNI0KMT_0_LC_12_12_5  (
            .in0(N__8766),
            .in1(N__8634),
            .in2(_gnd_net_),
            .in3(N__8581),
            .lcout(),
            .ltout(\uut.g1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.g0_2_LC_12_12_6 .C_ON=1'b0;
    defparam \uut.AR_BUF.g0_2_LC_12_12_6 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.g0_2_LC_12_12_6 .LUT_INIT=16'b1110101011000000;
    LogicCell40 \uut.AR_BUF.g0_2_LC_12_12_6  (
            .in0(N__7804),
            .in1(N__8597),
            .in2(N__7786),
            .in3(N__7782),
            .lcout(\uut.AR_BUF.g0_1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_RNIFFTC1_0_LC_12_12_7 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_RNIFFTC1_0_LC_12_12_7 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_RNIFFTC1_0_LC_12_12_7 .LUT_INIT=16'b1110000011000000;
    LogicCell40 \uut.seq.counter.T_1_RNIFFTC1_0_LC_12_12_7  (
            .in0(N__8765),
            .in1(N__8633),
            .in2(N__8601),
            .in3(N__8580),
            .lcout(\uut.program_counter_m_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.out_1_iv_0_LC_12_13_0 .C_ON=1'b0;
    defparam \uut.AR_BUF.out_1_iv_0_LC_12_13_0 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.out_1_iv_0_LC_12_13_0 .LUT_INIT=16'b1110111010101010;
    LogicCell40 \uut.AR_BUF.out_1_iv_0_LC_12_13_0  (
            .in0(N__8477),
            .in1(N__8430),
            .in2(_gnd_net_),
            .in3(N__8382),
            .lcout(),
            .ltout(\uut.AR_BUF.out_1_ivZ0Z_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.out_1_iv_2_1_LC_12_13_1 .C_ON=1'b0;
    defparam \uut.AR_BUF.out_1_iv_2_1_LC_12_13_1 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.out_1_iv_2_1_LC_12_13_1 .LUT_INIT=16'b1111111111111100;
    LogicCell40 \uut.AR_BUF.out_1_iv_2_1_LC_12_13_1  (
            .in0(_gnd_net_),
            .in1(N__9840),
            .in2(N__8308),
            .in3(N__8305),
            .lcout(),
            .ltout(\uut.out_1_iv_2_1_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.out_reg.ff4.q_LC_12_13_2 .C_ON=1'b0;
    defparam \uut.out_reg.ff4.q_LC_12_13_2 .SEQ_MODE=4'b1000;
    defparam \uut.out_reg.ff4.q_LC_12_13_2 .LUT_INIT=16'b1111110010101010;
    LogicCell40 \uut.out_reg.ff4.q_LC_12_13_2  (
            .in0(N__8157),
            .in1(N__8131),
            .in2(N__8290),
            .in3(N__8279),
            .lcout(LED4_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.out_reg.ff4.qC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mem.data_2_7_0__m15_LC_12_13_3 .C_ON=1'b0;
    defparam \uut.mem.data_2_7_0__m15_LC_12_13_3 .SEQ_MODE=4'b0000;
    defparam \uut.mem.data_2_7_0__m15_LC_12_13_3 .LUT_INIT=16'b0100100011001000;
    LogicCell40 \uut.mem.data_2_7_0__m15_LC_12_13_3  (
            .in0(N__9665),
            .in1(N__9535),
            .in2(N__9609),
            .in3(N__8845),
            .lcout(),
            .ltout(\uut.m15_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.AR_BUF.out_1_iv_3_LC_12_13_4 .C_ON=1'b0;
    defparam \uut.AR_BUF.out_1_iv_3_LC_12_13_4 .SEQ_MODE=4'b0000;
    defparam \uut.AR_BUF.out_1_iv_3_LC_12_13_4 .LUT_INIT=16'b1100110011001111;
    LogicCell40 \uut.AR_BUF.out_1_iv_3_LC_12_13_4  (
            .in0(_gnd_net_),
            .in1(N__8140),
            .in2(N__8134),
            .in3(N__8971),
            .lcout(\uut.out_1_iv_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mar.ff1.q_sbtinv_LC_12_13_5 .C_ON=1'b0;
    defparam \uut.mar.ff1.q_sbtinv_LC_12_13_5 .SEQ_MODE=4'b0000;
    defparam \uut.mar.ff1.q_sbtinv_LC_12_13_5 .LUT_INIT=16'b0000000011111111;
    LogicCell40 \uut.mar.ff1.q_sbtinv_LC_12_13_5  (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__8043),
            .lcout(\uut.mar.MAR_LD_0_1 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mar.ff3.q_LC_12_13_6 .C_ON=1'b0;
    defparam \uut.mar.ff3.q_LC_12_13_6 .SEQ_MODE=4'b1000;
    defparam \uut.mar.ff3.q_LC_12_13_6 .LUT_INIT=16'b1111111000001110;
    LogicCell40 \uut.mar.ff3.q_LC_12_13_6  (
            .in0(N__8121),
            .in1(N__8066),
            .in2(N__8047),
            .in3(N__9666),
            .lcout(\uut.mar_out_2 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.out_reg.ff4.qC_net ),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mem.data_2_7_0__g1_LC_12_13_7 .C_ON=1'b0;
    defparam \uut.mem.data_2_7_0__g1_LC_12_13_7 .SEQ_MODE=4'b0000;
    defparam \uut.mem.data_2_7_0__g1_LC_12_13_7 .LUT_INIT=16'b0110011011101110;
    LogicCell40 \uut.mem.data_2_7_0__g1_LC_12_13_7  (
            .in0(N__9590),
            .in1(N__9651),
            .in2(_gnd_net_),
            .in3(N__8844),
            .lcout(\uut.g1_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mar.ff4.q_ne_LC_12_14_0 .C_ON=1'b0;
    defparam \uut.mar.ff4.q_ne_LC_12_14_0 .SEQ_MODE=4'b1000;
    defparam \uut.mar.ff4.q_ne_LC_12_14_0 .LUT_INIT=16'b1111111111111110;
    LogicCell40 \uut.mar.ff4.q_ne_LC_12_14_0  (
            .in0(N__9851),
            .in1(N__9803),
            .in2(N__9772),
            .in3(N__9714),
            .lcout(\uut.mar_out_3 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.mar.ff4.q_neC_net ),
            .ce(N__8800),
            .sr(_gnd_net_));
    defparam \uut.mem.data_2_7_0__m6_LC_12_14_1 .C_ON=1'b0;
    defparam \uut.mem.data_2_7_0__m6_LC_12_14_1 .SEQ_MODE=4'b0000;
    defparam \uut.mem.data_2_7_0__m6_LC_12_14_1 .LUT_INIT=16'b0111111110100111;
    LogicCell40 \uut.mem.data_2_7_0__m6_LC_12_14_1  (
            .in0(N__9650),
            .in1(N__9571),
            .in2(N__9543),
            .in3(N__8827),
            .lcout(\uut.m6 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.seq.counter.T_1_fast_RNI38VD1_1_LC_12_14_2 .C_ON=1'b0;
    defparam \uut.seq.counter.T_1_fast_RNI38VD1_1_LC_12_14_2 .SEQ_MODE=4'b0000;
    defparam \uut.seq.counter.T_1_fast_RNI38VD1_1_LC_12_14_2 .LUT_INIT=16'b1000100010111011;
    LogicCell40 \uut.seq.counter.T_1_fast_RNI38VD1_1_LC_12_14_2  (
            .in0(N__9481),
            .in1(N__9464),
            .in2(_gnd_net_),
            .in3(N__9427),
            .lcout(\uut.un1_ROM_OE_0 ),
            .ltout(\uut.un1_ROM_OE_0_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mem.data_2_7_0__N_7_i_m_sx_LC_12_14_3 .C_ON=1'b0;
    defparam \uut.mem.data_2_7_0__N_7_i_m_sx_LC_12_14_3 .SEQ_MODE=4'b0000;
    defparam \uut.mem.data_2_7_0__N_7_i_m_sx_LC_12_14_3 .LUT_INIT=16'b1111111101010000;
    LogicCell40 \uut.mem.data_2_7_0__N_7_i_m_sx_LC_12_14_3  (
            .in0(N__9356),
            .in1(_gnd_net_),
            .in2(N__9313),
            .in3(N__9110),
            .lcout(),
            .ltout(\uut.mem.N_7_i_m_sx_cascade_ ),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mem.data_2_7_0__N_7_i_m_LC_12_14_4 .C_ON=1'b0;
    defparam \uut.mem.data_2_7_0__N_7_i_m_LC_12_14_4 .SEQ_MODE=4'b0000;
    defparam \uut.mem.data_2_7_0__N_7_i_m_LC_12_14_4 .LUT_INIT=16'b0000011100001111;
    LogicCell40 \uut.mem.data_2_7_0__N_7_i_m_LC_12_14_4  (
            .in0(N__9309),
            .in1(N__9298),
            .in2(N__9286),
            .in3(N__9283),
            .lcout(\uut.N_7_i_m ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam \uut.mar.ff1.q_ne_LC_12_14_5 .C_ON=1'b0;
    defparam \uut.mar.ff1.q_ne_LC_12_14_5 .SEQ_MODE=4'b1000;
    defparam \uut.mar.ff1.q_ne_LC_12_14_5 .LUT_INIT=16'b1110111011101111;
    LogicCell40 \uut.mar.ff1.q_ne_LC_12_14_5  (
            .in0(N__9241),
            .in1(N__9196),
            .in2(N__9133),
            .in3(N__8977),
            .lcout(\uut.mar_out_0 ),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(\INVuut.mar.ff4.q_neC_net ),
            .ce(N__8800),
            .sr(_gnd_net_));
endmodule // test
